magic
tech sky130A
magscale 1 2
timestamp 1746239859
<< checkpaint >>
rect -3932 -3932 23330 25474
<< viali >>
rect 2513 18921 2547 18955
rect 9689 18921 9723 18955
rect 2605 18853 2639 18887
rect 5273 18853 5307 18887
rect 8585 18853 8619 18887
rect 10793 18853 10827 18887
rect 1409 18717 1443 18751
rect 1777 18717 1811 18751
rect 2329 18717 2363 18751
rect 2789 18717 2823 18751
rect 2881 18717 2915 18751
rect 2973 18717 3007 18751
rect 3617 18717 3651 18751
rect 4169 18717 4203 18751
rect 4537 18717 4571 18751
rect 5089 18717 5123 18751
rect 5641 18717 5675 18751
rect 6561 18717 6595 18751
rect 6745 18717 6779 18751
rect 7297 18717 7331 18751
rect 7849 18717 7883 18751
rect 8401 18717 8435 18751
rect 8953 18717 8987 18751
rect 9505 18717 9539 18751
rect 10057 18717 10091 18751
rect 10609 18717 10643 18751
rect 11345 18717 11379 18751
rect 11897 18717 11931 18751
rect 12449 18717 12483 18751
rect 12817 18717 12851 18751
rect 13553 18717 13587 18751
rect 14289 18717 14323 18751
rect 14473 18717 14507 18751
rect 15025 18717 15059 18751
rect 15577 18717 15611 18751
rect 16313 18717 16347 18751
rect 16865 18717 16899 18751
rect 17233 18717 17267 18751
rect 17693 18717 17727 18751
rect 3157 18649 3191 18683
rect 1593 18581 1627 18615
rect 1961 18581 1995 18615
rect 3065 18581 3099 18615
rect 3433 18581 3467 18615
rect 3985 18581 4019 18615
rect 4721 18581 4755 18615
rect 5825 18581 5859 18615
rect 6377 18581 6411 18615
rect 6929 18581 6963 18615
rect 7481 18581 7515 18615
rect 8033 18581 8067 18615
rect 9137 18581 9171 18615
rect 10241 18581 10275 18615
rect 11161 18581 11195 18615
rect 11713 18581 11747 18615
rect 12265 18581 12299 18615
rect 13001 18581 13035 18615
rect 13369 18581 13403 18615
rect 14105 18581 14139 18615
rect 14657 18581 14691 18615
rect 15209 18581 15243 18615
rect 15761 18581 15795 18615
rect 16129 18581 16163 18615
rect 16681 18581 16715 18615
rect 17417 18581 17451 18615
rect 17877 18581 17911 18615
rect 3157 18377 3191 18411
rect 15117 18377 15151 18411
rect 3617 18309 3651 18343
rect 6653 18309 6687 18343
rect 11069 18309 11103 18343
rect 13001 18309 13035 18343
rect 13737 18309 13771 18343
rect 15761 18309 15795 18343
rect 1409 18241 1443 18275
rect 3433 18241 3467 18275
rect 3709 18241 3743 18275
rect 6377 18241 6411 18275
rect 8401 18241 8435 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 10701 18241 10735 18275
rect 10793 18241 10827 18275
rect 10885 18241 10919 18275
rect 12173 18241 12207 18275
rect 12725 18241 12759 18275
rect 12909 18241 12943 18275
rect 13185 18241 13219 18275
rect 13369 18241 13403 18275
rect 13461 18241 13495 18275
rect 13553 18241 13587 18275
rect 13829 18241 13863 18275
rect 15025 18241 15059 18275
rect 15301 18241 15335 18275
rect 15577 18241 15611 18275
rect 15853 18241 15887 18275
rect 15945 18241 15979 18275
rect 16129 18241 16163 18275
rect 16865 18241 16899 18275
rect 17877 18241 17911 18275
rect 1685 18173 1719 18207
rect 4077 18173 4111 18207
rect 4353 18173 4387 18207
rect 8677 18173 8711 18207
rect 10149 18173 10183 18207
rect 12265 18173 12299 18207
rect 12633 18173 12667 18207
rect 16037 18173 16071 18207
rect 16773 18173 16807 18207
rect 13645 18105 13679 18139
rect 17233 18105 17267 18139
rect 3249 18037 3283 18071
rect 5825 18037 5859 18071
rect 8125 18037 8159 18071
rect 10241 18037 10275 18071
rect 10793 18037 10827 18071
rect 11989 18037 12023 18071
rect 12817 18037 12851 18071
rect 15485 18037 15519 18071
rect 15669 18037 15703 18071
rect 17693 18037 17727 18071
rect 2421 17833 2455 17867
rect 6929 17833 6963 17867
rect 9505 17833 9539 17867
rect 13553 17833 13587 17867
rect 14105 17833 14139 17867
rect 5365 17765 5399 17799
rect 2697 17697 2731 17731
rect 3065 17697 3099 17731
rect 7113 17697 7147 17731
rect 8125 17697 8159 17731
rect 9689 17697 9723 17731
rect 11437 17697 11471 17731
rect 12081 17697 12115 17731
rect 15853 17697 15887 17731
rect 17877 17697 17911 17731
rect 2605 17629 2639 17663
rect 3157 17629 3191 17663
rect 3341 17629 3375 17663
rect 4997 17629 5031 17663
rect 5273 17629 5307 17663
rect 5365 17629 5399 17663
rect 5641 17629 5675 17663
rect 7205 17629 7239 17663
rect 7573 17629 7607 17663
rect 7665 17629 7699 17663
rect 7941 17629 7975 17663
rect 9781 17629 9815 17663
rect 10241 17629 10275 17663
rect 10425 17629 10459 17663
rect 11529 17629 11563 17663
rect 11805 17629 11839 17663
rect 5457 17561 5491 17595
rect 10149 17561 10183 17595
rect 15577 17561 15611 17595
rect 17601 17561 17635 17595
rect 3249 17493 3283 17527
rect 4813 17493 4847 17527
rect 5181 17493 5215 17527
rect 7757 17493 7791 17527
rect 10241 17493 10275 17527
rect 11161 17493 11195 17527
rect 16129 17493 16163 17527
rect 4445 17289 4479 17323
rect 7481 17289 7515 17323
rect 8401 17289 8435 17323
rect 15485 17289 15519 17323
rect 5089 17221 5123 17255
rect 7389 17221 7423 17255
rect 9873 17221 9907 17255
rect 14841 17221 14875 17255
rect 2789 17153 2823 17187
rect 4629 17153 4663 17187
rect 5181 17153 5215 17187
rect 5365 17153 5399 17187
rect 7297 17153 7331 17187
rect 7573 17153 7607 17187
rect 7665 17153 7699 17187
rect 7849 17153 7883 17187
rect 15301 17153 15335 17187
rect 2881 17085 2915 17119
rect 4721 17085 4755 17119
rect 10149 17085 10183 17119
rect 15209 17085 15243 17119
rect 3157 17017 3191 17051
rect 5273 16949 5307 16983
rect 7757 16949 7791 16983
rect 1409 16745 1443 16779
rect 16037 16745 16071 16779
rect 4353 16677 4387 16711
rect 7389 16677 7423 16711
rect 2881 16609 2915 16643
rect 3157 16609 3191 16643
rect 4813 16609 4847 16643
rect 5365 16609 5399 16643
rect 6837 16609 6871 16643
rect 7113 16609 7147 16643
rect 7665 16609 7699 16643
rect 9965 16609 9999 16643
rect 14289 16609 14323 16643
rect 17877 16609 17911 16643
rect 4721 16541 4755 16575
rect 7757 16541 7791 16575
rect 9873 16541 9907 16575
rect 12541 16541 12575 16575
rect 12633 16541 12667 16575
rect 12817 16473 12851 16507
rect 14565 16473 14599 16507
rect 17601 16473 17635 16507
rect 10241 16405 10275 16439
rect 12725 16405 12759 16439
rect 16129 16405 16163 16439
rect 14197 16201 14231 16235
rect 17249 16201 17283 16235
rect 4261 16133 4295 16167
rect 17049 16133 17083 16167
rect 4537 16065 4571 16099
rect 13369 16065 13403 16099
rect 13461 16065 13495 16099
rect 13645 16065 13679 16099
rect 14565 16065 14599 16099
rect 17509 16065 17543 16099
rect 11529 15997 11563 16031
rect 11805 15997 11839 16031
rect 13277 15997 13311 16031
rect 14657 15997 14691 16031
rect 17417 15929 17451 15963
rect 2789 15861 2823 15895
rect 13829 15861 13863 15895
rect 17233 15861 17267 15895
rect 17693 15861 17727 15895
rect 8309 15657 8343 15691
rect 12081 15657 12115 15691
rect 14749 15657 14783 15691
rect 16773 15589 16807 15623
rect 6561 15521 6595 15555
rect 10241 15521 10275 15555
rect 11989 15521 12023 15555
rect 12357 15521 12391 15555
rect 13093 15521 13127 15555
rect 13553 15521 13587 15555
rect 1777 15453 1811 15487
rect 5181 15453 5215 15487
rect 5273 15453 5307 15487
rect 5641 15453 5675 15487
rect 5825 15453 5859 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 12265 15453 12299 15487
rect 12725 15453 12759 15487
rect 13001 15453 13035 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 14657 15453 14691 15487
rect 14841 15453 14875 15487
rect 16773 15453 16807 15487
rect 17049 15453 17083 15487
rect 17141 15453 17175 15487
rect 17325 15453 17359 15487
rect 5457 15385 5491 15419
rect 6837 15385 6871 15419
rect 10517 15385 10551 15419
rect 1961 15317 1995 15351
rect 5365 15317 5399 15351
rect 5825 15317 5859 15351
rect 9229 15317 9263 15351
rect 13369 15317 13403 15351
rect 16957 15317 16991 15351
rect 17233 15317 17267 15351
rect 5641 15113 5675 15147
rect 6929 15113 6963 15147
rect 10057 15113 10091 15147
rect 10425 15113 10459 15147
rect 15025 15113 15059 15147
rect 15669 15113 15703 15147
rect 10793 15045 10827 15079
rect 15761 15045 15795 15079
rect 3893 14977 3927 15011
rect 5917 14977 5951 15011
rect 6101 14977 6135 15011
rect 6193 14977 6227 15011
rect 6561 14977 6595 15011
rect 8217 14977 8251 15011
rect 10241 14977 10275 15011
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 10885 14977 10919 15011
rect 11805 14977 11839 15011
rect 14657 14977 14691 15011
rect 15301 14977 15335 15011
rect 15485 14977 15519 15011
rect 15577 14977 15611 15011
rect 15669 14977 15703 15011
rect 15945 14977 15979 15011
rect 1409 14909 1443 14943
rect 1685 14909 1719 14943
rect 4169 14909 4203 14943
rect 6469 14909 6503 14943
rect 8493 14909 8527 14943
rect 9965 14909 9999 14943
rect 14565 14909 14599 14943
rect 15117 14841 15151 14875
rect 3157 14773 3191 14807
rect 5733 14773 5767 14807
rect 10701 14773 10735 14807
rect 14381 14773 14415 14807
rect 2053 14569 2087 14603
rect 7297 14569 7331 14603
rect 8953 14569 8987 14603
rect 15853 14569 15887 14603
rect 2237 14433 2271 14467
rect 2973 14433 3007 14467
rect 9137 14433 9171 14467
rect 9597 14433 9631 14467
rect 14105 14433 14139 14467
rect 17693 14433 17727 14467
rect 2329 14365 2363 14399
rect 3157 14365 3191 14399
rect 3433 14365 3467 14399
rect 4353 14365 4387 14399
rect 4629 14365 4663 14399
rect 9229 14365 9263 14399
rect 6377 14297 6411 14331
rect 8769 14297 8803 14331
rect 11805 14297 11839 14331
rect 13553 14297 13587 14331
rect 14381 14297 14415 14331
rect 15945 14297 15979 14331
rect 2697 14229 2731 14263
rect 3341 14229 3375 14263
rect 2881 14025 2915 14059
rect 5089 14025 5123 14059
rect 5733 14025 5767 14059
rect 6377 14025 6411 14059
rect 3157 13957 3191 13991
rect 11161 13957 11195 13991
rect 11805 13957 11839 13991
rect 15025 13957 15059 13991
rect 16865 13957 16899 13991
rect 17049 13957 17083 13991
rect 2513 13889 2547 13923
rect 2697 13889 2731 13923
rect 2881 13889 2915 13923
rect 2973 13889 3007 13923
rect 5273 13889 5307 13923
rect 8125 13889 8159 13923
rect 11069 13889 11103 13923
rect 11345 13889 11379 13923
rect 11713 13889 11747 13923
rect 11989 13889 12023 13923
rect 16773 13889 16807 13923
rect 17141 13889 17175 13923
rect 17325 13889 17359 13923
rect 5365 13821 5399 13855
rect 7849 13821 7883 13855
rect 17233 13821 17267 13855
rect 2605 13685 2639 13719
rect 11253 13685 11287 13719
rect 12173 13685 12207 13719
rect 16957 13685 16991 13719
rect 10149 13481 10183 13515
rect 12817 13481 12851 13515
rect 2513 13345 2547 13379
rect 7021 13345 7055 13379
rect 8769 13345 8803 13379
rect 9229 13345 9263 13379
rect 12173 13345 12207 13379
rect 13001 13345 13035 13379
rect 17601 13345 17635 13379
rect 17877 13345 17911 13379
rect 2421 13277 2455 13311
rect 4813 13277 4847 13311
rect 4905 13277 4939 13311
rect 9321 13277 9355 13311
rect 11897 13277 11931 13311
rect 12265 13277 12299 13311
rect 13093 13277 13127 13311
rect 5089 13209 5123 13243
rect 7297 13209 7331 13243
rect 11621 13209 11655 13243
rect 11989 13209 12023 13243
rect 2053 13141 2087 13175
rect 4997 13141 5031 13175
rect 8953 13141 8987 13175
rect 12633 13141 12667 13175
rect 16129 13141 16163 13175
rect 5733 12937 5767 12971
rect 6929 12937 6963 12971
rect 12173 12937 12207 12971
rect 12817 12937 12851 12971
rect 17417 12937 17451 12971
rect 1685 12869 1719 12903
rect 9229 12869 9263 12903
rect 1409 12801 1443 12835
rect 3249 12801 3283 12835
rect 5273 12801 5307 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 6561 12801 6595 12835
rect 8953 12801 8987 12835
rect 11989 12801 12023 12835
rect 12173 12801 12207 12835
rect 14565 12801 14599 12835
rect 16405 12801 16439 12835
rect 16865 12801 16899 12835
rect 17601 12801 17635 12835
rect 17785 12801 17819 12835
rect 17877 12801 17911 12835
rect 3525 12733 3559 12767
rect 5089 12733 5123 12767
rect 5365 12733 5399 12767
rect 5917 12733 5951 12767
rect 6469 12733 6503 12767
rect 14289 12733 14323 12767
rect 14657 12733 14691 12767
rect 16129 12733 16163 12767
rect 16957 12733 16991 12767
rect 17325 12733 17359 12767
rect 3157 12597 3191 12631
rect 4997 12597 5031 12631
rect 10701 12597 10735 12631
rect 16681 12597 16715 12631
rect 5549 12393 5583 12427
rect 10425 12393 10459 12427
rect 17509 12393 17543 12427
rect 15761 12257 15795 12291
rect 5089 12189 5123 12223
rect 5365 12189 5399 12223
rect 7941 12189 7975 12223
rect 8217 12189 8251 12223
rect 8401 12189 8435 12223
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 10241 12189 10275 12223
rect 10333 12189 10367 12223
rect 10609 12189 10643 12223
rect 10885 12189 10919 12223
rect 12633 12189 12667 12223
rect 12909 12189 12943 12223
rect 3249 12121 3283 12155
rect 10517 12121 10551 12155
rect 12725 12121 12759 12155
rect 16037 12121 16071 12155
rect 3525 12053 3559 12087
rect 5181 12053 5215 12087
rect 8033 12053 8067 12087
rect 8493 12053 8527 12087
rect 10701 12053 10735 12087
rect 11069 12053 11103 12087
rect 13093 12053 13127 12087
rect 8125 11849 8159 11883
rect 8861 11849 8895 11883
rect 9045 11849 9079 11883
rect 13553 11849 13587 11883
rect 14749 11849 14783 11883
rect 2513 11781 2547 11815
rect 8953 11781 8987 11815
rect 2421 11713 2455 11747
rect 2697 11713 2731 11747
rect 3341 11713 3375 11747
rect 6377 11713 6411 11747
rect 8401 11713 8435 11747
rect 9137 11713 9171 11747
rect 9229 11713 9263 11747
rect 11345 11713 11379 11747
rect 11805 11713 11839 11747
rect 14381 11713 14415 11747
rect 3433 11645 3467 11679
rect 6653 11645 6687 11679
rect 8217 11645 8251 11679
rect 8493 11645 8527 11679
rect 12081 11645 12115 11679
rect 14473 11645 14507 11679
rect 3709 11577 3743 11611
rect 2605 11509 2639 11543
rect 9873 11509 9907 11543
rect 3433 11305 3467 11339
rect 4997 11305 5031 11339
rect 11161 11305 11195 11339
rect 12265 11305 12299 11339
rect 14749 11305 14783 11339
rect 7941 11237 7975 11271
rect 13185 11237 13219 11271
rect 2237 11169 2271 11203
rect 3249 11169 3283 11203
rect 6469 11169 6503 11203
rect 6745 11169 6779 11203
rect 8401 11169 8435 11203
rect 12449 11169 12483 11203
rect 16773 11169 16807 11203
rect 2329 11101 2363 11135
rect 2697 11101 2731 11135
rect 2789 11101 2823 11135
rect 3065 11101 3099 11135
rect 3341 11101 3375 11135
rect 3525 11101 3559 11135
rect 8309 11101 8343 11135
rect 9413 11101 9447 11135
rect 11253 11101 11287 11135
rect 11437 11101 11471 11135
rect 12541 11101 12575 11135
rect 12909 11101 12943 11135
rect 13001 11101 13035 11135
rect 13369 11101 13403 11135
rect 13553 11101 13587 11135
rect 14657 11101 14691 11135
rect 14841 11101 14875 11135
rect 16681 11101 16715 11135
rect 9689 11033 9723 11067
rect 13093 11033 13127 11067
rect 13277 11033 13311 11067
rect 2053 10965 2087 10999
rect 2881 10965 2915 10999
rect 11253 10965 11287 10999
rect 13369 10965 13403 10999
rect 16313 10965 16347 10999
rect 3157 10761 3191 10795
rect 9965 10761 9999 10795
rect 10609 10761 10643 10795
rect 15025 10761 15059 10795
rect 15669 10761 15703 10795
rect 1685 10693 1719 10727
rect 4077 10693 4111 10727
rect 6469 10693 6503 10727
rect 15485 10693 15519 10727
rect 15761 10693 15795 10727
rect 17141 10693 17175 10727
rect 10149 10625 10183 10659
rect 10241 10625 10275 10659
rect 14565 10625 14599 10659
rect 15117 10625 15151 10659
rect 15301 10625 15335 10659
rect 15577 10625 15611 10659
rect 15669 10625 15703 10659
rect 15945 10625 15979 10659
rect 16773 10625 16807 10659
rect 1409 10557 1443 10591
rect 3801 10557 3835 10591
rect 6745 10557 6779 10591
rect 14657 10557 14691 10591
rect 5549 10421 5583 10455
rect 14381 10421 14415 10455
rect 15853 10217 15887 10251
rect 6561 10149 6595 10183
rect 10517 10081 10551 10115
rect 12541 10081 12575 10115
rect 14381 10081 14415 10115
rect 16405 10081 16439 10115
rect 4629 10013 4663 10047
rect 4721 10013 4755 10047
rect 4905 10013 4939 10047
rect 6285 10013 6319 10047
rect 6837 10013 6871 10047
rect 10425 10013 10459 10047
rect 12449 10013 12483 10047
rect 14105 10013 14139 10047
rect 16129 10013 16163 10047
rect 7205 9945 7239 9979
rect 5089 9877 5123 9911
rect 10793 9877 10827 9911
rect 12817 9877 12851 9911
rect 17877 9877 17911 9911
rect 5457 9673 5491 9707
rect 6929 9673 6963 9707
rect 13277 9673 13311 9707
rect 2421 9605 2455 9639
rect 7481 9605 7515 9639
rect 10057 9605 10091 9639
rect 11805 9605 11839 9639
rect 16773 9605 16807 9639
rect 17325 9605 17359 9639
rect 2329 9537 2363 9571
rect 2605 9537 2639 9571
rect 6561 9537 6595 9571
rect 9965 9537 9999 9571
rect 10241 9537 10275 9571
rect 17233 9537 17267 9571
rect 17509 9537 17543 9571
rect 3709 9469 3743 9503
rect 3985 9469 4019 9503
rect 6653 9469 6687 9503
rect 7205 9469 7239 9503
rect 8953 9469 8987 9503
rect 11529 9469 11563 9503
rect 2329 9333 2363 9367
rect 10149 9333 10183 9367
rect 17049 9333 17083 9367
rect 17693 9333 17727 9367
rect 7205 9129 7239 9163
rect 10701 9129 10735 9163
rect 15853 9129 15887 9163
rect 8033 9061 8067 9095
rect 3157 8993 3191 9027
rect 6377 8993 6411 9027
rect 6561 8993 6595 9027
rect 7389 8993 7423 9027
rect 8953 8993 8987 9027
rect 13921 8993 13955 9027
rect 14105 8993 14139 9027
rect 16497 8993 16531 9027
rect 1409 8925 1443 8959
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 6101 8925 6135 8959
rect 6285 8925 6319 8959
rect 6653 8925 6687 8959
rect 7113 8925 7147 8959
rect 7297 8925 7331 8959
rect 7573 8925 7607 8959
rect 7849 8925 7883 8959
rect 7941 8925 7975 8959
rect 8217 8925 8251 8959
rect 10977 8925 11011 8959
rect 11253 8925 11287 8959
rect 16589 8925 16623 8959
rect 17049 8925 17083 8959
rect 1685 8857 1719 8891
rect 6009 8857 6043 8891
rect 8125 8857 8159 8891
rect 9229 8857 9263 8891
rect 13645 8857 13679 8891
rect 14381 8857 14415 8891
rect 17141 8857 17175 8891
rect 17325 8857 17359 8891
rect 6101 8789 6135 8823
rect 7021 8789 7055 8823
rect 7757 8789 7791 8823
rect 10793 8789 10827 8823
rect 11161 8789 11195 8823
rect 12173 8789 12207 8823
rect 16313 8789 16347 8823
rect 16957 8789 16991 8823
rect 17049 8789 17083 8823
rect 2881 8585 2915 8619
rect 4169 8585 4203 8619
rect 5089 8585 5123 8619
rect 9873 8585 9907 8619
rect 10517 8585 10551 8619
rect 12633 8585 12667 8619
rect 15945 8585 15979 8619
rect 5181 8517 5215 8551
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 4353 8449 4387 8483
rect 4905 8449 4939 8483
rect 4997 8449 5031 8483
rect 10057 8449 10091 8483
rect 10609 8449 10643 8483
rect 10793 8449 10827 8483
rect 12541 8449 12575 8483
rect 12817 8449 12851 8483
rect 14473 8449 14507 8483
rect 14657 8449 14691 8483
rect 16681 8449 16715 8483
rect 16865 8449 16899 8483
rect 4445 8381 4479 8415
rect 4813 8381 4847 8415
rect 10149 8381 10183 8415
rect 2513 8245 2547 8279
rect 10701 8245 10735 8279
rect 13001 8245 13035 8279
rect 16773 8245 16807 8279
rect 1685 8041 1719 8075
rect 6929 8041 6963 8075
rect 12449 8041 12483 8075
rect 14197 8041 14231 8075
rect 17509 8041 17543 8075
rect 2329 7905 2363 7939
rect 4353 7905 4387 7939
rect 5181 7905 5215 7939
rect 14565 7905 14599 7939
rect 15761 7905 15795 7939
rect 16037 7905 16071 7939
rect 1869 7837 1903 7871
rect 1961 7837 1995 7871
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 4261 7837 4295 7871
rect 8769 7837 8803 7871
rect 13921 7837 13955 7871
rect 14473 7837 14507 7871
rect 5457 7769 5491 7803
rect 2513 7701 2547 7735
rect 4629 7701 4663 7735
rect 7481 7701 7515 7735
rect 9781 7497 9815 7531
rect 15025 7497 15059 7531
rect 5273 7429 5307 7463
rect 5549 7361 5583 7395
rect 9321 7361 9355 7395
rect 9597 7361 9631 7395
rect 9873 7361 9907 7395
rect 10333 7361 10367 7395
rect 12541 7361 12575 7395
rect 14749 7361 14783 7395
rect 14933 7361 14967 7395
rect 15025 7361 15059 7395
rect 15209 7361 15243 7395
rect 17049 7361 17083 7395
rect 1961 7293 1995 7327
rect 2237 7293 2271 7327
rect 9045 7293 9079 7327
rect 10425 7293 10459 7327
rect 16957 7293 16991 7327
rect 3801 7225 3835 7259
rect 3709 7157 3743 7191
rect 7573 7157 7607 7191
rect 9413 7157 9447 7191
rect 10057 7157 10091 7191
rect 14841 7157 14875 7191
rect 16773 7157 16807 7191
rect 9597 6953 9631 6987
rect 10136 6953 10170 6987
rect 13829 6953 13863 6987
rect 15853 6953 15887 6987
rect 16392 6953 16426 6987
rect 2053 6885 2087 6919
rect 1777 6817 1811 6851
rect 5273 6817 5307 6851
rect 7021 6817 7055 6851
rect 9413 6817 9447 6851
rect 9873 6817 9907 6851
rect 11713 6817 11747 6851
rect 13461 6817 13495 6851
rect 14565 6817 14599 6851
rect 14933 6817 14967 6851
rect 16129 6817 16163 6851
rect 1685 6749 1719 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 8493 6749 8527 6783
rect 8769 6749 8803 6783
rect 9321 6749 9355 6783
rect 13553 6749 13587 6783
rect 13737 6749 13771 6783
rect 13829 6749 13863 6783
rect 14473 6749 14507 6783
rect 15209 6749 15243 6783
rect 15393 6749 15427 6783
rect 15669 6749 15703 6783
rect 16037 6749 16071 6783
rect 5549 6681 5583 6715
rect 8585 6681 8619 6715
rect 11989 6681 12023 6715
rect 15761 6681 15795 6715
rect 15945 6681 15979 6715
rect 8401 6613 8435 6647
rect 8677 6613 8711 6647
rect 8953 6613 8987 6647
rect 11621 6613 11655 6647
rect 14289 6613 14323 6647
rect 15577 6613 15611 6647
rect 17877 6613 17911 6647
rect 11989 6409 12023 6443
rect 12633 6409 12667 6443
rect 15485 6409 15519 6443
rect 14013 6341 14047 6375
rect 2973 6273 3007 6307
rect 3065 6273 3099 6307
rect 3525 6273 3559 6307
rect 3709 6273 3743 6307
rect 12173 6273 12207 6307
rect 13737 6273 13771 6307
rect 3433 6205 3467 6239
rect 12265 6205 12299 6239
rect 2789 6069 2823 6103
rect 3617 6069 3651 6103
rect 3801 5865 3835 5899
rect 5549 5865 5583 5899
rect 7849 5797 7883 5831
rect 1685 5729 1719 5763
rect 1961 5729 1995 5763
rect 5365 5729 5399 5763
rect 6837 5729 6871 5763
rect 9229 5729 9263 5763
rect 12357 5729 12391 5763
rect 16037 5729 16071 5763
rect 1593 5661 1627 5695
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 5273 5661 5307 5695
rect 6745 5661 6779 5695
rect 6929 5661 6963 5695
rect 7389 5661 7423 5695
rect 7573 5661 7607 5695
rect 7665 5661 7699 5695
rect 7941 5661 7975 5695
rect 8033 5661 8067 5695
rect 9321 5661 9355 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 10977 5661 11011 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 12265 5661 12299 5695
rect 15945 5661 15979 5695
rect 16497 5661 16531 5695
rect 16589 5661 16623 5695
rect 7205 5593 7239 5627
rect 7757 5593 7791 5627
rect 11345 5593 11379 5627
rect 16773 5593 16807 5627
rect 1409 5525 1443 5559
rect 3433 5525 3467 5559
rect 4169 5525 4203 5559
rect 8953 5525 8987 5559
rect 11161 5525 11195 5559
rect 11437 5525 11471 5559
rect 12633 5525 12667 5559
rect 15761 5525 15795 5559
rect 16405 5525 16439 5559
rect 16681 5525 16715 5559
rect 7021 5321 7055 5355
rect 9321 5321 9355 5355
rect 11161 5321 11195 5355
rect 14197 5321 14231 5355
rect 16129 5321 16163 5355
rect 16497 5321 16531 5355
rect 3525 5253 3559 5287
rect 5917 5253 5951 5287
rect 13829 5253 13863 5287
rect 3157 5185 3191 5219
rect 3249 5185 3283 5219
rect 3341 5185 3375 5219
rect 3985 5185 4019 5219
rect 6193 5185 6227 5219
rect 7573 5185 7607 5219
rect 9413 5185 9447 5219
rect 11897 5185 11931 5219
rect 15945 5185 15979 5219
rect 16037 5185 16071 5219
rect 16313 5185 16347 5219
rect 17233 5185 17267 5219
rect 1409 5117 1443 5151
rect 2881 5117 2915 5151
rect 3893 5117 3927 5151
rect 6561 5117 6595 5151
rect 6653 5117 6687 5151
rect 7849 5117 7883 5151
rect 9689 5117 9723 5151
rect 11805 5117 11839 5151
rect 12357 5117 12391 5151
rect 14105 5117 14139 5151
rect 15669 5117 15703 5151
rect 17141 5117 17175 5151
rect 3433 5049 3467 5083
rect 3617 5049 3651 5083
rect 11529 5049 11563 5083
rect 16865 5049 16899 5083
rect 4445 4981 4479 5015
rect 6377 4981 6411 5015
rect 7849 4777 7883 4811
rect 10517 4777 10551 4811
rect 11345 4777 11379 4811
rect 16681 4777 16715 4811
rect 16865 4777 16899 4811
rect 6101 4641 6135 4675
rect 6377 4641 6411 4675
rect 10701 4641 10735 4675
rect 11161 4641 11195 4675
rect 14933 4641 14967 4675
rect 10793 4573 10827 4607
rect 11253 4573 11287 4607
rect 11437 4573 11471 4607
rect 16773 4573 16807 4607
rect 16957 4573 16991 4607
rect 15209 4505 15243 4539
rect 15117 2465 15151 2499
rect 14565 2397 14599 2431
<< metal1 >>
rect 1104 19066 18216 19088
rect 1104 19014 1918 19066
rect 1970 19014 1982 19066
rect 2034 19014 2046 19066
rect 2098 19014 2110 19066
rect 2162 19014 2174 19066
rect 2226 19014 2238 19066
rect 2290 19014 7918 19066
rect 7970 19014 7982 19066
rect 8034 19014 8046 19066
rect 8098 19014 8110 19066
rect 8162 19014 8174 19066
rect 8226 19014 8238 19066
rect 8290 19014 13918 19066
rect 13970 19014 13982 19066
rect 14034 19014 14046 19066
rect 14098 19014 14110 19066
rect 14162 19014 14174 19066
rect 14226 19014 14238 19066
rect 14290 19014 18216 19066
rect 1104 18992 18216 19014
rect 2501 18955 2559 18961
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 4430 18952 4436 18964
rect 2547 18924 4436 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 4430 18912 4436 18924
rect 4488 18912 4494 18964
rect 9677 18955 9735 18961
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 12434 18952 12440 18964
rect 9723 18924 12440 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 1578 18844 1584 18896
rect 1636 18884 1642 18896
rect 2593 18887 2651 18893
rect 2593 18884 2605 18887
rect 1636 18856 2605 18884
rect 1636 18844 1642 18856
rect 2593 18853 2605 18856
rect 2639 18853 2651 18887
rect 2593 18847 2651 18853
rect 5261 18887 5319 18893
rect 5261 18853 5273 18887
rect 5307 18884 5319 18887
rect 6822 18884 6828 18896
rect 5307 18856 6828 18884
rect 5307 18853 5319 18856
rect 5261 18847 5319 18853
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 8573 18887 8631 18893
rect 8573 18853 8585 18887
rect 8619 18884 8631 18887
rect 9398 18884 9404 18896
rect 8619 18856 9404 18884
rect 8619 18853 8631 18856
rect 8573 18847 8631 18853
rect 9398 18844 9404 18856
rect 9456 18844 9462 18896
rect 10781 18887 10839 18893
rect 10781 18853 10793 18887
rect 10827 18884 10839 18887
rect 12618 18884 12624 18896
rect 10827 18856 12624 18884
rect 10827 18853 10839 18856
rect 10781 18847 10839 18853
rect 12618 18844 12624 18856
rect 12676 18844 12682 18896
rect 5350 18816 5356 18828
rect 2884 18788 5356 18816
rect 1118 18708 1124 18760
rect 1176 18748 1182 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 1176 18720 1409 18748
rect 1176 18708 1182 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1670 18708 1676 18760
rect 1728 18748 1734 18760
rect 1765 18751 1823 18757
rect 1765 18748 1777 18751
rect 1728 18720 1777 18748
rect 1728 18708 1734 18720
rect 1765 18717 1777 18720
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 2314 18708 2320 18760
rect 2372 18708 2378 18760
rect 2774 18708 2780 18760
rect 2832 18708 2838 18760
rect 2884 18757 2912 18788
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 2869 18751 2927 18757
rect 2869 18717 2881 18751
rect 2915 18717 2927 18751
rect 2869 18711 2927 18717
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18748 3019 18751
rect 3007 18720 3280 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 3142 18640 3148 18692
rect 3200 18640 3206 18692
rect 3252 18680 3280 18720
rect 3326 18708 3332 18760
rect 3384 18748 3390 18760
rect 3605 18751 3663 18757
rect 3605 18748 3617 18751
rect 3384 18720 3617 18748
rect 3384 18708 3390 18720
rect 3605 18717 3617 18720
rect 3651 18717 3663 18751
rect 3605 18711 3663 18717
rect 3878 18708 3884 18760
rect 3936 18748 3942 18760
rect 4157 18751 4215 18757
rect 4157 18748 4169 18751
rect 3936 18720 4169 18748
rect 3936 18708 3942 18720
rect 4157 18717 4169 18720
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 4522 18708 4528 18760
rect 4580 18708 4586 18760
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 5077 18751 5135 18757
rect 5077 18748 5089 18751
rect 5040 18720 5089 18748
rect 5040 18708 5046 18720
rect 5077 18717 5089 18720
rect 5123 18717 5135 18751
rect 5077 18711 5135 18717
rect 5626 18708 5632 18760
rect 5684 18708 5690 18760
rect 6086 18708 6092 18760
rect 6144 18748 6150 18760
rect 6549 18751 6607 18757
rect 6549 18748 6561 18751
rect 6144 18720 6561 18748
rect 6144 18708 6150 18720
rect 6549 18717 6561 18720
rect 6595 18717 6607 18751
rect 6549 18711 6607 18717
rect 6638 18708 6644 18760
rect 6696 18748 6702 18760
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6696 18720 6745 18748
rect 6696 18708 6702 18720
rect 6733 18717 6745 18720
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 7282 18708 7288 18760
rect 7340 18708 7346 18760
rect 7834 18708 7840 18760
rect 7892 18708 7898 18760
rect 8386 18708 8392 18760
rect 8444 18708 8450 18760
rect 8938 18708 8944 18760
rect 8996 18708 9002 18760
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 10042 18708 10048 18760
rect 10100 18708 10106 18760
rect 10502 18708 10508 18760
rect 10560 18748 10566 18760
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10560 18720 10609 18748
rect 10560 18708 10566 18720
rect 10597 18717 10609 18720
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 11112 18720 11345 18748
rect 11112 18708 11118 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11664 18720 11897 18748
rect 11664 18708 11670 18720
rect 11885 18717 11897 18720
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12437 18751 12495 18757
rect 12437 18748 12449 18751
rect 12216 18720 12449 18748
rect 12216 18708 12222 18720
rect 12437 18717 12449 18720
rect 12483 18717 12495 18751
rect 12437 18711 12495 18717
rect 12710 18708 12716 18760
rect 12768 18748 12774 18760
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12768 18720 12817 18748
rect 12768 18708 12774 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 13538 18708 13544 18760
rect 13596 18708 13602 18760
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13872 18720 14289 18748
rect 13872 18708 13878 18720
rect 14277 18717 14289 18720
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 14458 18708 14464 18760
rect 14516 18708 14522 18760
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 15562 18708 15568 18760
rect 15620 18708 15626 18760
rect 16298 18708 16304 18760
rect 16356 18708 16362 18760
rect 16850 18708 16856 18760
rect 16908 18708 16914 18760
rect 17218 18708 17224 18760
rect 17276 18708 17282 18760
rect 17678 18708 17684 18760
rect 17736 18708 17742 18760
rect 10686 18680 10692 18692
rect 3252 18652 3740 18680
rect 3712 18624 3740 18652
rect 9140 18652 10692 18680
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 1581 18615 1639 18621
rect 1581 18612 1593 18615
rect 1544 18584 1593 18612
rect 1544 18572 1550 18584
rect 1581 18581 1593 18584
rect 1627 18581 1639 18615
rect 1581 18575 1639 18581
rect 1762 18572 1768 18624
rect 1820 18612 1826 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1820 18584 1961 18612
rect 1820 18572 1826 18584
rect 1949 18581 1961 18584
rect 1995 18581 2007 18615
rect 1949 18575 2007 18581
rect 3050 18572 3056 18624
rect 3108 18572 3114 18624
rect 3418 18572 3424 18624
rect 3476 18572 3482 18624
rect 3694 18572 3700 18624
rect 3752 18612 3758 18624
rect 3973 18615 4031 18621
rect 3973 18612 3985 18615
rect 3752 18584 3985 18612
rect 3752 18572 3758 18584
rect 3973 18581 3985 18584
rect 4019 18581 4031 18615
rect 3973 18575 4031 18581
rect 4709 18615 4767 18621
rect 4709 18581 4721 18615
rect 4755 18612 4767 18615
rect 5166 18612 5172 18624
rect 4755 18584 5172 18612
rect 4755 18581 4767 18584
rect 4709 18575 4767 18581
rect 5166 18572 5172 18584
rect 5224 18572 5230 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 5813 18615 5871 18621
rect 5813 18612 5825 18615
rect 5592 18584 5825 18612
rect 5592 18572 5598 18584
rect 5813 18581 5825 18584
rect 5859 18581 5871 18615
rect 5813 18575 5871 18581
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 6365 18615 6423 18621
rect 6365 18612 6377 18615
rect 5960 18584 6377 18612
rect 5960 18572 5966 18584
rect 6365 18581 6377 18584
rect 6411 18581 6423 18615
rect 6365 18575 6423 18581
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7098 18612 7104 18624
rect 6963 18584 7104 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 7466 18572 7472 18624
rect 7524 18572 7530 18624
rect 7650 18572 7656 18624
rect 7708 18612 7714 18624
rect 9140 18621 9168 18652
rect 10686 18640 10692 18652
rect 10744 18640 10750 18692
rect 8021 18615 8079 18621
rect 8021 18612 8033 18615
rect 7708 18584 8033 18612
rect 7708 18572 7714 18584
rect 8021 18581 8033 18584
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 9125 18615 9183 18621
rect 9125 18581 9137 18615
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10229 18615 10287 18621
rect 10229 18612 10241 18615
rect 10192 18584 10241 18612
rect 10192 18572 10198 18584
rect 10229 18581 10241 18584
rect 10275 18581 10287 18615
rect 10229 18575 10287 18581
rect 11149 18615 11207 18621
rect 11149 18581 11161 18615
rect 11195 18612 11207 18615
rect 11330 18612 11336 18624
rect 11195 18584 11336 18612
rect 11195 18581 11207 18584
rect 11149 18575 11207 18581
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 12253 18615 12311 18621
rect 12253 18612 12265 18615
rect 12216 18584 12265 18612
rect 12216 18572 12222 18584
rect 12253 18581 12265 18584
rect 12299 18581 12311 18615
rect 12253 18575 12311 18581
rect 12986 18572 12992 18624
rect 13044 18572 13050 18624
rect 13354 18572 13360 18624
rect 13412 18572 13418 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 13780 18584 14105 18612
rect 13780 18572 13786 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 14608 18584 14657 18612
rect 14608 18572 14614 18584
rect 14645 18581 14657 18584
rect 14691 18581 14703 18615
rect 14645 18575 14703 18581
rect 15197 18615 15255 18621
rect 15197 18581 15209 18615
rect 15243 18612 15255 18615
rect 15562 18612 15568 18624
rect 15243 18584 15568 18612
rect 15243 18581 15255 18584
rect 15197 18575 15255 18581
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15746 18572 15752 18624
rect 15804 18572 15810 18624
rect 15838 18572 15844 18624
rect 15896 18612 15902 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15896 18584 16129 18612
rect 15896 18572 15902 18584
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 16117 18575 16175 18581
rect 16666 18572 16672 18624
rect 16724 18572 16730 18624
rect 17310 18572 17316 18624
rect 17368 18612 17374 18624
rect 17405 18615 17463 18621
rect 17405 18612 17417 18615
rect 17368 18584 17417 18612
rect 17368 18572 17374 18584
rect 17405 18581 17417 18584
rect 17451 18581 17463 18615
rect 17405 18575 17463 18581
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 17865 18615 17923 18621
rect 17865 18612 17877 18615
rect 17828 18584 17877 18612
rect 17828 18572 17834 18584
rect 17865 18581 17877 18584
rect 17911 18581 17923 18615
rect 17865 18575 17923 18581
rect 1104 18522 18216 18544
rect 1104 18470 2658 18522
rect 2710 18470 2722 18522
rect 2774 18470 2786 18522
rect 2838 18470 2850 18522
rect 2902 18470 2914 18522
rect 2966 18470 2978 18522
rect 3030 18470 8658 18522
rect 8710 18470 8722 18522
rect 8774 18470 8786 18522
rect 8838 18470 8850 18522
rect 8902 18470 8914 18522
rect 8966 18470 8978 18522
rect 9030 18470 14658 18522
rect 14710 18470 14722 18522
rect 14774 18470 14786 18522
rect 14838 18470 14850 18522
rect 14902 18470 14914 18522
rect 14966 18470 14978 18522
rect 15030 18470 18216 18522
rect 1104 18448 18216 18470
rect 3142 18368 3148 18420
rect 3200 18368 3206 18420
rect 7282 18408 7288 18420
rect 4724 18380 6316 18408
rect 2406 18300 2412 18352
rect 2464 18300 2470 18352
rect 1397 18275 1455 18281
rect 1397 18241 1409 18275
rect 1443 18241 1455 18275
rect 3160 18272 3188 18368
rect 3605 18343 3663 18349
rect 3605 18309 3617 18343
rect 3651 18340 3663 18343
rect 3786 18340 3792 18352
rect 3651 18312 3792 18340
rect 3651 18309 3663 18312
rect 3605 18303 3663 18309
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 4724 18340 4752 18380
rect 3988 18312 4830 18340
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 3160 18244 3433 18272
rect 1397 18235 1455 18241
rect 3421 18241 3433 18244
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 1412 18068 1440 18235
rect 3694 18232 3700 18284
rect 3752 18232 3758 18284
rect 1670 18164 1676 18216
rect 1728 18164 1734 18216
rect 2406 18164 2412 18216
rect 2464 18204 2470 18216
rect 3988 18204 4016 18312
rect 2464 18176 4016 18204
rect 4065 18207 4123 18213
rect 2464 18164 2470 18176
rect 4065 18173 4077 18207
rect 4111 18173 4123 18207
rect 4065 18167 4123 18173
rect 3142 18136 3148 18148
rect 2746 18108 3148 18136
rect 2746 18068 2774 18108
rect 3142 18096 3148 18108
rect 3200 18136 3206 18148
rect 4080 18136 4108 18167
rect 4338 18164 4344 18216
rect 4396 18164 4402 18216
rect 6288 18204 6316 18380
rect 6380 18380 7288 18408
rect 6380 18281 6408 18380
rect 7282 18368 7288 18380
rect 7340 18408 7346 18420
rect 8202 18408 8208 18420
rect 7340 18380 8208 18408
rect 7340 18368 7346 18380
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 13354 18408 13360 18420
rect 8312 18380 8800 18408
rect 6641 18343 6699 18349
rect 6641 18309 6653 18343
rect 6687 18340 6699 18343
rect 6914 18340 6920 18352
rect 6687 18312 6920 18340
rect 6687 18309 6699 18312
rect 6641 18303 6699 18309
rect 6914 18300 6920 18312
rect 6972 18300 6978 18352
rect 6365 18275 6423 18281
rect 6365 18241 6377 18275
rect 6411 18241 6423 18275
rect 8312 18272 8340 18380
rect 8772 18340 8800 18380
rect 11072 18380 13360 18408
rect 9122 18340 9128 18352
rect 8772 18312 9128 18340
rect 9122 18300 9128 18312
rect 9180 18300 9186 18352
rect 11072 18349 11100 18380
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 13446 18368 13452 18420
rect 13504 18408 13510 18420
rect 15105 18411 15163 18417
rect 15105 18408 15117 18411
rect 13504 18380 15117 18408
rect 13504 18368 13510 18380
rect 15105 18377 15117 18380
rect 15151 18377 15163 18411
rect 15105 18371 15163 18377
rect 11057 18343 11115 18349
rect 11057 18340 11069 18343
rect 10704 18312 11069 18340
rect 7774 18258 8340 18272
rect 6365 18235 6423 18241
rect 7760 18244 8340 18258
rect 8389 18275 8447 18281
rect 7760 18204 7788 18244
rect 8389 18241 8401 18275
rect 8435 18241 8447 18275
rect 8389 18235 8447 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 6288 18176 7788 18204
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8404 18204 8432 18235
rect 8260 18176 8432 18204
rect 8260 18164 8266 18176
rect 8662 18164 8668 18216
rect 8720 18164 8726 18216
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18204 10195 18207
rect 10428 18204 10456 18235
rect 10594 18232 10600 18284
rect 10652 18232 10658 18284
rect 10704 18281 10732 18312
rect 11057 18309 11069 18312
rect 11103 18309 11115 18343
rect 12989 18343 13047 18349
rect 12989 18340 13001 18343
rect 11057 18303 11115 18309
rect 12728 18312 13001 18340
rect 12728 18281 12756 18312
rect 12989 18309 13001 18312
rect 13035 18309 13047 18343
rect 13722 18340 13728 18352
rect 12989 18303 13047 18309
rect 13464 18312 13728 18340
rect 10689 18275 10747 18281
rect 10689 18241 10701 18275
rect 10735 18241 10747 18275
rect 10689 18235 10747 18241
rect 10781 18275 10839 18281
rect 10781 18241 10793 18275
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 12161 18275 12219 18281
rect 12161 18241 12173 18275
rect 12207 18272 12219 18275
rect 12713 18275 12771 18281
rect 12713 18272 12725 18275
rect 12207 18244 12725 18272
rect 12207 18241 12219 18244
rect 12161 18235 12219 18241
rect 12713 18241 12725 18244
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 10796 18204 10824 18235
rect 10183 18176 10824 18204
rect 10183 18173 10195 18176
rect 10137 18167 10195 18173
rect 3200 18108 4108 18136
rect 3200 18096 3206 18108
rect 10594 18096 10600 18148
rect 10652 18136 10658 18148
rect 10888 18136 10916 18235
rect 12250 18164 12256 18216
rect 12308 18164 12314 18216
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18204 12679 18207
rect 12912 18204 12940 18235
rect 12667 18176 12940 18204
rect 13188 18204 13216 18235
rect 13354 18232 13360 18284
rect 13412 18232 13418 18284
rect 13464 18281 13492 18312
rect 13722 18300 13728 18312
rect 13780 18300 13786 18352
rect 15749 18343 15807 18349
rect 15749 18340 15761 18343
rect 15028 18312 15761 18340
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 13538 18232 13544 18284
rect 13596 18232 13602 18284
rect 13817 18275 13875 18281
rect 13817 18241 13829 18275
rect 13863 18241 13875 18275
rect 13817 18235 13875 18241
rect 13556 18204 13584 18232
rect 13188 18176 13584 18204
rect 13832 18204 13860 18235
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 15028 18281 15056 18312
rect 15749 18309 15761 18312
rect 15795 18309 15807 18343
rect 15749 18303 15807 18309
rect 15013 18275 15071 18281
rect 15013 18272 15025 18275
rect 14608 18244 15025 18272
rect 14608 18232 14614 18244
rect 15013 18241 15025 18244
rect 15059 18241 15071 18275
rect 15013 18235 15071 18241
rect 15194 18232 15200 18284
rect 15252 18272 15258 18284
rect 15289 18275 15347 18281
rect 15565 18278 15623 18281
rect 15289 18272 15301 18275
rect 15252 18244 15301 18272
rect 15252 18232 15258 18244
rect 15289 18241 15301 18244
rect 15335 18272 15347 18275
rect 15488 18275 15623 18278
rect 15488 18272 15577 18275
rect 15335 18250 15577 18272
rect 15335 18244 15516 18250
rect 15335 18241 15347 18244
rect 15289 18235 15347 18241
rect 15565 18241 15577 18250
rect 15611 18241 15623 18275
rect 15841 18275 15899 18281
rect 15841 18272 15853 18275
rect 15565 18235 15623 18241
rect 15672 18244 15853 18272
rect 15378 18204 15384 18216
rect 13832 18176 15384 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 10652 18108 10916 18136
rect 12912 18136 12940 18176
rect 15378 18164 15384 18176
rect 15436 18204 15442 18216
rect 15672 18204 15700 18244
rect 15841 18241 15853 18244
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 15930 18232 15936 18284
rect 15988 18232 15994 18284
rect 16114 18232 16120 18284
rect 16172 18232 16178 18284
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16264 18244 16865 18272
rect 16264 18232 16270 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 18230 18272 18236 18284
rect 17911 18244 18236 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 18230 18232 18236 18244
rect 18288 18232 18294 18284
rect 15436 18176 15700 18204
rect 16025 18207 16083 18213
rect 15436 18164 15442 18176
rect 16025 18173 16037 18207
rect 16071 18204 16083 18207
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 16071 18176 16773 18204
rect 16071 18173 16083 18176
rect 16025 18167 16083 18173
rect 16761 18173 16773 18176
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 12912 18108 13645 18136
rect 10652 18096 10658 18108
rect 13633 18105 13645 18108
rect 13679 18105 13691 18139
rect 16114 18136 16120 18148
rect 13633 18099 13691 18105
rect 15488 18108 16120 18136
rect 1412 18040 2774 18068
rect 3234 18028 3240 18080
rect 3292 18028 3298 18080
rect 5810 18028 5816 18080
rect 5868 18028 5874 18080
rect 7834 18028 7840 18080
rect 7892 18068 7898 18080
rect 8113 18071 8171 18077
rect 8113 18068 8125 18071
rect 7892 18040 8125 18068
rect 7892 18028 7898 18040
rect 8113 18037 8125 18040
rect 8159 18037 8171 18071
rect 8113 18031 8171 18037
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 10468 18040 10793 18068
rect 10468 18028 10474 18040
rect 10781 18037 10793 18040
rect 10827 18037 10839 18071
rect 10781 18031 10839 18037
rect 11977 18071 12035 18077
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12066 18068 12072 18080
rect 12023 18040 12072 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 12802 18028 12808 18080
rect 12860 18028 12866 18080
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 15488 18077 15516 18108
rect 16114 18096 16120 18108
rect 16172 18096 16178 18148
rect 17221 18139 17279 18145
rect 17221 18105 17233 18139
rect 17267 18136 17279 18139
rect 17586 18136 17592 18148
rect 17267 18108 17592 18136
rect 17267 18105 17279 18108
rect 17221 18099 17279 18105
rect 17586 18096 17592 18108
rect 17644 18096 17650 18148
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 15344 18040 15485 18068
rect 15344 18028 15350 18040
rect 15473 18037 15485 18040
rect 15519 18037 15531 18071
rect 15473 18031 15531 18037
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 15930 18068 15936 18080
rect 15712 18040 15936 18068
rect 15712 18028 15718 18040
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 17678 18028 17684 18080
rect 17736 18028 17742 18080
rect 1104 17978 18216 18000
rect 1104 17926 1918 17978
rect 1970 17926 1982 17978
rect 2034 17926 2046 17978
rect 2098 17926 2110 17978
rect 2162 17926 2174 17978
rect 2226 17926 2238 17978
rect 2290 17926 7918 17978
rect 7970 17926 7982 17978
rect 8034 17926 8046 17978
rect 8098 17926 8110 17978
rect 8162 17926 8174 17978
rect 8226 17926 8238 17978
rect 8290 17926 13918 17978
rect 13970 17926 13982 17978
rect 14034 17926 14046 17978
rect 14098 17926 14110 17978
rect 14162 17926 14174 17978
rect 14226 17926 14238 17978
rect 14290 17926 18216 17978
rect 1104 17904 18216 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2409 17867 2467 17873
rect 2409 17864 2421 17867
rect 1728 17836 2421 17864
rect 1728 17824 1734 17836
rect 2409 17833 2421 17836
rect 2455 17833 2467 17867
rect 2409 17827 2467 17833
rect 6914 17824 6920 17876
rect 6972 17824 6978 17876
rect 8662 17824 8668 17876
rect 8720 17864 8726 17876
rect 9493 17867 9551 17873
rect 9493 17864 9505 17867
rect 8720 17836 9505 17864
rect 8720 17824 8726 17836
rect 9493 17833 9505 17836
rect 9539 17833 9551 17867
rect 12802 17864 12808 17876
rect 9493 17827 9551 17833
rect 11440 17836 12808 17864
rect 5258 17756 5264 17808
rect 5316 17796 5322 17808
rect 5353 17799 5411 17805
rect 5353 17796 5365 17799
rect 5316 17768 5365 17796
rect 5316 17756 5322 17768
rect 5353 17765 5365 17768
rect 5399 17765 5411 17799
rect 5353 17759 5411 17765
rect 2498 17688 2504 17740
rect 2556 17728 2562 17740
rect 2685 17731 2743 17737
rect 2685 17728 2697 17731
rect 2556 17700 2697 17728
rect 2556 17688 2562 17700
rect 2685 17697 2697 17700
rect 2731 17697 2743 17731
rect 2685 17691 2743 17697
rect 3050 17688 3056 17740
rect 3108 17728 3114 17740
rect 7101 17731 7159 17737
rect 3108 17700 3188 17728
rect 3108 17688 3114 17700
rect 3160 17669 3188 17700
rect 5000 17700 5672 17728
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17629 2651 17663
rect 2593 17623 2651 17629
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17629 3203 17663
rect 3145 17623 3203 17629
rect 2608 17592 2636 17623
rect 3234 17620 3240 17672
rect 3292 17660 3298 17672
rect 5000 17669 5028 17700
rect 3329 17663 3387 17669
rect 3329 17660 3341 17663
rect 3292 17632 3341 17660
rect 3292 17620 3298 17632
rect 3329 17629 3341 17632
rect 3375 17629 3387 17663
rect 3329 17623 3387 17629
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17629 5043 17663
rect 4985 17623 5043 17629
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 5261 17663 5319 17669
rect 5261 17660 5273 17663
rect 5224 17632 5273 17660
rect 5224 17620 5230 17632
rect 5261 17629 5273 17632
rect 5307 17629 5319 17663
rect 5261 17623 5319 17629
rect 3252 17592 3280 17620
rect 2608 17564 3280 17592
rect 3786 17552 3792 17604
rect 3844 17592 3850 17604
rect 5276 17592 5304 17623
rect 5350 17620 5356 17672
rect 5408 17620 5414 17672
rect 5644 17669 5672 17700
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7742 17728 7748 17740
rect 7147 17700 7748 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 7742 17688 7748 17700
rect 7800 17728 7806 17740
rect 11440 17737 11468 17836
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 13538 17824 13544 17876
rect 13596 17824 13602 17876
rect 14093 17867 14151 17873
rect 14093 17833 14105 17867
rect 14139 17864 14151 17867
rect 15194 17864 15200 17876
rect 14139 17836 15200 17864
rect 14139 17833 14151 17836
rect 14093 17827 14151 17833
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 8113 17731 8171 17737
rect 8113 17728 8125 17731
rect 7800 17700 8125 17728
rect 7800 17688 7806 17700
rect 8113 17697 8125 17700
rect 8159 17697 8171 17731
rect 8113 17691 8171 17697
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 11425 17731 11483 17737
rect 9723 17700 10272 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 10244 17672 10272 17700
rect 11425 17697 11437 17731
rect 11471 17697 11483 17731
rect 11425 17691 11483 17697
rect 12066 17688 12072 17740
rect 12124 17688 12130 17740
rect 14550 17688 14556 17740
rect 14608 17728 14614 17740
rect 15841 17731 15899 17737
rect 15841 17728 15853 17731
rect 14608 17700 15853 17728
rect 14608 17688 14614 17700
rect 15841 17697 15853 17700
rect 15887 17728 15899 17731
rect 17862 17728 17868 17740
rect 15887 17700 17868 17728
rect 15887 17697 15899 17700
rect 15841 17691 15899 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 5810 17660 5816 17672
rect 5675 17632 5816 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 5810 17620 5816 17632
rect 5868 17620 5874 17672
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 7558 17620 7564 17672
rect 7616 17620 7622 17672
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 5445 17595 5503 17601
rect 5445 17592 5457 17595
rect 3844 17564 5212 17592
rect 5276 17564 5457 17592
rect 3844 17552 3850 17564
rect 3234 17484 3240 17536
rect 3292 17484 3298 17536
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 5184 17533 5212 17564
rect 5445 17561 5457 17564
rect 5491 17561 5503 17595
rect 5445 17555 5503 17561
rect 6822 17552 6828 17604
rect 6880 17592 6886 17604
rect 7668 17592 7696 17623
rect 7834 17620 7840 17672
rect 7892 17660 7898 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7892 17632 7941 17660
rect 7892 17620 7898 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 9766 17620 9772 17672
rect 9824 17620 9830 17672
rect 10226 17620 10232 17672
rect 10284 17620 10290 17672
rect 10410 17620 10416 17672
rect 10468 17620 10474 17672
rect 11517 17663 11575 17669
rect 11517 17629 11529 17663
rect 11563 17629 11575 17663
rect 11517 17623 11575 17629
rect 6880 17564 7696 17592
rect 10137 17595 10195 17601
rect 6880 17552 6886 17564
rect 10137 17561 10149 17595
rect 10183 17592 10195 17595
rect 10428 17592 10456 17620
rect 10183 17564 10456 17592
rect 11532 17592 11560 17623
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11664 17632 11805 17660
rect 11664 17620 11670 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 13814 17592 13820 17604
rect 11532 17564 12296 17592
rect 13294 17564 13820 17592
rect 10183 17561 10195 17564
rect 10137 17555 10195 17561
rect 12268 17536 12296 17564
rect 13814 17552 13820 17564
rect 13872 17592 13878 17604
rect 13872 17564 14398 17592
rect 13872 17552 13878 17564
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 15565 17595 15623 17601
rect 15565 17592 15577 17595
rect 15528 17564 15577 17592
rect 15528 17552 15534 17564
rect 15565 17561 15577 17564
rect 15611 17561 15623 17595
rect 15565 17555 15623 17561
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 16356 17564 16422 17592
rect 16356 17552 16362 17564
rect 17586 17552 17592 17604
rect 17644 17552 17650 17604
rect 4801 17527 4859 17533
rect 4801 17524 4813 17527
rect 4672 17496 4813 17524
rect 4672 17484 4678 17496
rect 4801 17493 4813 17496
rect 4847 17493 4859 17527
rect 4801 17487 4859 17493
rect 5169 17527 5227 17533
rect 5169 17493 5181 17527
rect 5215 17524 5227 17527
rect 7745 17527 7803 17533
rect 7745 17524 7757 17527
rect 5215 17496 7757 17524
rect 5215 17493 5227 17496
rect 5169 17487 5227 17493
rect 7745 17493 7757 17496
rect 7791 17493 7803 17527
rect 7745 17487 7803 17493
rect 10226 17484 10232 17536
rect 10284 17484 10290 17536
rect 11146 17484 11152 17536
rect 11204 17484 11210 17536
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 16117 17527 16175 17533
rect 16117 17524 16129 17527
rect 12308 17496 16129 17524
rect 12308 17484 12314 17496
rect 16117 17493 16129 17496
rect 16163 17493 16175 17527
rect 16117 17487 16175 17493
rect 1104 17434 18216 17456
rect 1104 17382 2658 17434
rect 2710 17382 2722 17434
rect 2774 17382 2786 17434
rect 2838 17382 2850 17434
rect 2902 17382 2914 17434
rect 2966 17382 2978 17434
rect 3030 17382 8658 17434
rect 8710 17382 8722 17434
rect 8774 17382 8786 17434
rect 8838 17382 8850 17434
rect 8902 17382 8914 17434
rect 8966 17382 8978 17434
rect 9030 17382 14658 17434
rect 14710 17382 14722 17434
rect 14774 17382 14786 17434
rect 14838 17382 14850 17434
rect 14902 17382 14914 17434
rect 14966 17382 14978 17434
rect 15030 17382 18216 17434
rect 1104 17360 18216 17382
rect 4338 17280 4344 17332
rect 4396 17320 4402 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 4396 17292 4445 17320
rect 4396 17280 4402 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 4433 17283 4491 17289
rect 7469 17323 7527 17329
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 7558 17320 7564 17332
rect 7515 17292 7564 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 8389 17323 8447 17329
rect 8389 17289 8401 17323
rect 8435 17320 8447 17323
rect 9766 17320 9772 17332
rect 8435 17292 9772 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 15470 17280 15476 17332
rect 15528 17280 15534 17332
rect 5077 17255 5135 17261
rect 5077 17221 5089 17255
rect 5123 17252 5135 17255
rect 5123 17224 5304 17252
rect 5123 17221 5135 17224
rect 5077 17215 5135 17221
rect 5276 17196 5304 17224
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 7377 17255 7435 17261
rect 7377 17252 7389 17255
rect 6880 17224 7389 17252
rect 6880 17212 6886 17224
rect 7377 17221 7389 17224
rect 7423 17221 7435 17255
rect 7576 17252 7604 17280
rect 7576 17224 7696 17252
rect 7377 17215 7435 17221
rect 1394 17144 1400 17196
rect 1452 17184 1458 17196
rect 2498 17184 2504 17196
rect 1452 17156 2504 17184
rect 1452 17144 1458 17156
rect 2498 17144 2504 17156
rect 2556 17184 2562 17196
rect 2777 17187 2835 17193
rect 2777 17184 2789 17187
rect 2556 17156 2789 17184
rect 2556 17144 2562 17156
rect 2777 17153 2789 17156
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 5169 17187 5227 17193
rect 5169 17184 5181 17187
rect 4672 17156 5181 17184
rect 4672 17144 4678 17156
rect 5169 17153 5181 17156
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 7668 17193 7696 17224
rect 7742 17212 7748 17264
rect 7800 17252 7806 17264
rect 7800 17224 7880 17252
rect 7800 17212 7806 17224
rect 7852 17193 7880 17224
rect 9122 17212 9128 17264
rect 9180 17212 9186 17264
rect 9861 17255 9919 17261
rect 9861 17221 9873 17255
rect 9907 17252 9919 17255
rect 11146 17252 11152 17264
rect 9907 17224 11152 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 11146 17212 11152 17224
rect 11204 17212 11210 17264
rect 14829 17255 14887 17261
rect 14829 17221 14841 17255
rect 14875 17252 14887 17255
rect 15654 17252 15660 17264
rect 14875 17224 15660 17252
rect 14875 17221 14887 17224
rect 14829 17215 14887 17221
rect 15654 17212 15660 17224
rect 15712 17212 15718 17264
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5316 17156 5365 17184
rect 5316 17144 5322 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17153 7711 17187
rect 7653 17147 7711 17153
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 3234 17116 3240 17128
rect 2915 17088 3240 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 4706 17076 4712 17128
rect 4764 17076 4770 17128
rect 3145 17051 3203 17057
rect 3145 17017 3157 17051
rect 3191 17048 3203 17051
rect 4246 17048 4252 17060
rect 3191 17020 4252 17048
rect 3191 17017 3203 17020
rect 3145 17011 3203 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 7300 17048 7328 17147
rect 7576 17116 7604 17147
rect 15286 17144 15292 17196
rect 15344 17144 15350 17196
rect 7742 17116 7748 17128
rect 7576 17088 7748 17116
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 11514 17116 11520 17128
rect 10183 17088 11520 17116
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 15197 17119 15255 17125
rect 15197 17085 15209 17119
rect 15243 17116 15255 17119
rect 16206 17116 16212 17128
rect 15243 17088 16212 17116
rect 15243 17085 15255 17088
rect 15197 17079 15255 17085
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 7300 17020 8892 17048
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 5261 16983 5319 16989
rect 5261 16980 5273 16983
rect 4856 16952 5273 16980
rect 4856 16940 4862 16952
rect 5261 16949 5273 16952
rect 5307 16949 5319 16983
rect 5261 16943 5319 16949
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 7745 16983 7803 16989
rect 7745 16980 7757 16983
rect 7708 16952 7757 16980
rect 7708 16940 7714 16952
rect 7745 16949 7757 16952
rect 7791 16949 7803 16983
rect 8864 16980 8892 17020
rect 10870 16980 10876 16992
rect 8864 16952 10876 16980
rect 7745 16943 7803 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 1104 16890 18216 16912
rect 1104 16838 1918 16890
rect 1970 16838 1982 16890
rect 2034 16838 2046 16890
rect 2098 16838 2110 16890
rect 2162 16838 2174 16890
rect 2226 16838 2238 16890
rect 2290 16838 7918 16890
rect 7970 16838 7982 16890
rect 8034 16838 8046 16890
rect 8098 16838 8110 16890
rect 8162 16838 8174 16890
rect 8226 16838 8238 16890
rect 8290 16838 13918 16890
rect 13970 16838 13982 16890
rect 14034 16838 14046 16890
rect 14098 16838 14110 16890
rect 14162 16838 14174 16890
rect 14226 16838 14238 16890
rect 14290 16838 18216 16890
rect 1104 16816 18216 16838
rect 1394 16736 1400 16788
rect 1452 16736 1458 16788
rect 16025 16779 16083 16785
rect 16025 16745 16037 16779
rect 16071 16776 16083 16779
rect 16206 16776 16212 16788
rect 16071 16748 16212 16776
rect 16071 16745 16083 16748
rect 16025 16739 16083 16745
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 4341 16711 4399 16717
rect 4341 16708 4353 16711
rect 3068 16680 4353 16708
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16640 2927 16643
rect 3068 16640 3096 16680
rect 4341 16677 4353 16680
rect 4387 16677 4399 16711
rect 7377 16711 7435 16717
rect 7377 16708 7389 16711
rect 4341 16671 4399 16677
rect 7024 16680 7389 16708
rect 2915 16612 3096 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 3142 16600 3148 16652
rect 3200 16600 3206 16652
rect 4798 16600 4804 16652
rect 4856 16600 4862 16652
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16640 6883 16643
rect 7024 16640 7052 16680
rect 7377 16677 7389 16680
rect 7423 16677 7435 16711
rect 7377 16671 7435 16677
rect 6871 16612 7052 16640
rect 7101 16643 7159 16649
rect 6871 16609 6883 16612
rect 6825 16603 6883 16609
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 7282 16640 7288 16652
rect 7147 16612 7288 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 4706 16532 4712 16584
rect 4764 16572 4770 16584
rect 5368 16572 5396 16603
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 7650 16600 7656 16652
rect 7708 16600 7714 16652
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10226 16640 10232 16652
rect 9999 16612 10232 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 14277 16643 14335 16649
rect 10928 16612 11008 16640
rect 10928 16600 10934 16612
rect 4764 16544 5396 16572
rect 4764 16532 4770 16544
rect 7190 16532 7196 16584
rect 7248 16572 7254 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7248 16544 7757 16572
rect 7248 16532 7254 16544
rect 7745 16541 7757 16544
rect 7791 16572 7803 16575
rect 7834 16572 7840 16584
rect 7791 16544 7840 16572
rect 7791 16541 7803 16544
rect 7745 16535 7803 16541
rect 7834 16532 7840 16544
rect 7892 16532 7898 16584
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9824 16544 9873 16572
rect 9824 16532 9830 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 10980 16572 11008 16612
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14550 16640 14556 16652
rect 14323 16612 14556 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 17862 16600 17868 16652
rect 17920 16600 17926 16652
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 10980 16544 12541 16572
rect 9861 16535 9919 16541
rect 12529 16541 12541 16544
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 13078 16572 13084 16584
rect 12667 16544 13084 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 2406 16464 2412 16516
rect 2464 16504 2470 16516
rect 4062 16504 4068 16516
rect 2464 16476 4068 16504
rect 2464 16464 2470 16476
rect 4062 16464 4068 16476
rect 4120 16504 4126 16516
rect 12805 16507 12863 16513
rect 4120 16476 5658 16504
rect 4120 16464 4126 16476
rect 12805 16473 12817 16507
rect 12851 16504 12863 16507
rect 13262 16504 13268 16516
rect 12851 16476 13268 16504
rect 12851 16473 12863 16476
rect 12805 16467 12863 16473
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 14182 16464 14188 16516
rect 14240 16504 14246 16516
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 14240 16476 14565 16504
rect 14240 16464 14246 16476
rect 14553 16473 14565 16476
rect 14599 16473 14611 16507
rect 16298 16504 16304 16516
rect 14553 16467 14611 16473
rect 14752 16476 15042 16504
rect 16040 16476 16304 16504
rect 10229 16439 10287 16445
rect 10229 16405 10241 16439
rect 10275 16436 10287 16439
rect 10502 16436 10508 16448
rect 10275 16408 10508 16436
rect 10275 16405 10287 16408
rect 10229 16399 10287 16405
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 12710 16396 12716 16448
rect 12768 16396 12774 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14752 16436 14780 16476
rect 15286 16436 15292 16448
rect 13872 16408 15292 16436
rect 13872 16396 13878 16408
rect 15286 16396 15292 16408
rect 15344 16436 15350 16448
rect 16040 16436 16068 16476
rect 16298 16464 16304 16476
rect 16356 16504 16362 16516
rect 16356 16476 16422 16504
rect 16356 16464 16362 16476
rect 17586 16464 17592 16516
rect 17644 16464 17650 16516
rect 15344 16408 16068 16436
rect 15344 16396 15350 16408
rect 16114 16396 16120 16448
rect 16172 16396 16178 16448
rect 1104 16346 18216 16368
rect 1104 16294 2658 16346
rect 2710 16294 2722 16346
rect 2774 16294 2786 16346
rect 2838 16294 2850 16346
rect 2902 16294 2914 16346
rect 2966 16294 2978 16346
rect 3030 16294 8658 16346
rect 8710 16294 8722 16346
rect 8774 16294 8786 16346
rect 8838 16294 8850 16346
rect 8902 16294 8914 16346
rect 8966 16294 8978 16346
rect 9030 16294 14658 16346
rect 14710 16294 14722 16346
rect 14774 16294 14786 16346
rect 14838 16294 14850 16346
rect 14902 16294 14914 16346
rect 14966 16294 14978 16346
rect 15030 16294 18216 16346
rect 1104 16272 18216 16294
rect 4062 16192 4068 16244
rect 4120 16192 4126 16244
rect 13814 16232 13820 16244
rect 12176 16204 13820 16232
rect 4080 16164 4108 16192
rect 3818 16136 4108 16164
rect 4246 16124 4252 16176
rect 4304 16124 4310 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 12176 16164 12204 16204
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 14182 16192 14188 16244
rect 14240 16192 14246 16244
rect 16114 16192 16120 16244
rect 16172 16232 16178 16244
rect 17237 16235 17295 16241
rect 17237 16232 17249 16235
rect 16172 16204 17249 16232
rect 16172 16192 16178 16204
rect 17237 16201 17249 16204
rect 17283 16201 17295 16235
rect 17237 16195 17295 16201
rect 11112 16136 12282 16164
rect 11112 16124 11118 16136
rect 13262 16124 13268 16176
rect 13320 16164 13326 16176
rect 13320 16136 13676 16164
rect 13320 16124 13326 16136
rect 4525 16099 4583 16105
rect 4525 16065 4537 16099
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 3234 15988 3240 16040
rect 3292 16028 3298 16040
rect 3878 16028 3884 16040
rect 3292 16000 3884 16028
rect 3292 15988 3298 16000
rect 3878 15988 3884 16000
rect 3936 16028 3942 16040
rect 4540 16028 4568 16059
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13136 16068 13369 16096
rect 13136 16056 13142 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13446 16056 13452 16108
rect 13504 16096 13510 16108
rect 13648 16105 13676 16136
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 16816 16136 17049 16164
rect 16816 16124 16822 16136
rect 17037 16133 17049 16136
rect 17083 16133 17095 16167
rect 17678 16164 17684 16176
rect 17037 16127 17095 16133
rect 17328 16136 17684 16164
rect 13633 16099 13691 16105
rect 13504 16068 13584 16096
rect 13504 16056 13510 16068
rect 3936 16000 4568 16028
rect 3936 15988 3942 16000
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 11793 16031 11851 16037
rect 11572 16000 11652 16028
rect 11572 15988 11578 16000
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 2777 15895 2835 15901
rect 2777 15892 2789 15895
rect 2372 15864 2789 15892
rect 2372 15852 2378 15864
rect 2777 15861 2789 15864
rect 2823 15861 2835 15895
rect 11624 15892 11652 16000
rect 11793 15997 11805 16031
rect 11839 16028 11851 16031
rect 11882 16028 11888 16040
rect 11839 16000 11888 16028
rect 11839 15997 11851 16000
rect 11793 15991 11851 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 13262 15988 13268 16040
rect 13320 15988 13326 16040
rect 13556 15960 13584 16068
rect 13633 16065 13645 16099
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16096 14611 16099
rect 15102 16096 15108 16108
rect 14599 16068 15108 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 16028 14703 16031
rect 14734 16028 14740 16040
rect 14691 16000 14740 16028
rect 14691 15997 14703 16000
rect 14645 15991 14703 15997
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 15470 15960 15476 15972
rect 13556 15932 15476 15960
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 17328 15960 17356 16136
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 17497 16099 17555 16105
rect 17497 16096 17509 16099
rect 17420 16068 17509 16096
rect 17420 15969 17448 16068
rect 17497 16065 17509 16068
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 17236 15932 17356 15960
rect 17405 15963 17463 15969
rect 11790 15892 11796 15904
rect 11624 15864 11796 15892
rect 2777 15855 2835 15861
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 13688 15864 13829 15892
rect 13688 15852 13694 15864
rect 13817 15861 13829 15864
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 17236 15901 17264 15932
rect 17405 15929 17417 15963
rect 17451 15929 17463 15963
rect 17405 15923 17463 15929
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 17092 15864 17233 15892
rect 17092 15852 17098 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 17586 15892 17592 15904
rect 17368 15864 17592 15892
rect 17368 15852 17374 15864
rect 17586 15852 17592 15864
rect 17644 15892 17650 15904
rect 17681 15895 17739 15901
rect 17681 15892 17693 15895
rect 17644 15864 17693 15892
rect 17644 15852 17650 15864
rect 17681 15861 17693 15864
rect 17727 15861 17739 15895
rect 17681 15855 17739 15861
rect 1104 15802 18216 15824
rect 1104 15750 1918 15802
rect 1970 15750 1982 15802
rect 2034 15750 2046 15802
rect 2098 15750 2110 15802
rect 2162 15750 2174 15802
rect 2226 15750 2238 15802
rect 2290 15750 7918 15802
rect 7970 15750 7982 15802
rect 8034 15750 8046 15802
rect 8098 15750 8110 15802
rect 8162 15750 8174 15802
rect 8226 15750 8238 15802
rect 8290 15750 13918 15802
rect 13970 15750 13982 15802
rect 14034 15750 14046 15802
rect 14098 15750 14110 15802
rect 14162 15750 14174 15802
rect 14226 15750 14238 15802
rect 14290 15750 18216 15802
rect 1104 15728 18216 15750
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 7892 15660 8309 15688
rect 7892 15648 7898 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 8297 15651 8355 15657
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 12069 15691 12127 15697
rect 12069 15688 12081 15691
rect 11940 15660 12081 15688
rect 11940 15648 11946 15660
rect 12069 15657 12081 15660
rect 12115 15657 12127 15691
rect 12069 15651 12127 15657
rect 14734 15648 14740 15700
rect 14792 15648 14798 15700
rect 12710 15580 12716 15632
rect 12768 15620 12774 15632
rect 13446 15620 13452 15632
rect 12768 15592 13452 15620
rect 12768 15580 12774 15592
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 16761 15623 16819 15629
rect 16761 15589 16773 15623
rect 16807 15589 16819 15623
rect 16761 15583 16819 15589
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 6178 15552 6184 15564
rect 5592 15524 6184 15552
rect 5592 15512 5598 15524
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15552 6607 15555
rect 7282 15552 7288 15564
rect 6595 15524 7288 15552
rect 6595 15521 6607 15524
rect 6549 15515 6607 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 10229 15555 10287 15561
rect 9048 15524 9904 15552
rect 934 15444 940 15496
rect 992 15484 998 15496
rect 1765 15487 1823 15493
rect 1765 15484 1777 15487
rect 992 15456 1777 15484
rect 992 15444 998 15456
rect 1765 15453 1777 15456
rect 1811 15453 1823 15487
rect 1765 15447 1823 15453
rect 4798 15444 4804 15496
rect 4856 15484 4862 15496
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 4856 15456 5181 15484
rect 4856 15444 4862 15456
rect 5169 15453 5181 15456
rect 5215 15453 5227 15487
rect 5169 15447 5227 15453
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15484 5319 15487
rect 5552 15484 5580 15512
rect 5307 15456 5580 15484
rect 5629 15487 5687 15493
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 5629 15453 5641 15487
rect 5675 15453 5687 15487
rect 5629 15447 5687 15453
rect 5445 15419 5503 15425
rect 5445 15385 5457 15419
rect 5491 15416 5503 15419
rect 5534 15416 5540 15428
rect 5491 15388 5540 15416
rect 5491 15385 5503 15388
rect 5445 15379 5503 15385
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 5644 15416 5672 15447
rect 5718 15444 5724 15496
rect 5776 15484 5782 15496
rect 5813 15487 5871 15493
rect 5813 15484 5825 15487
rect 5776 15456 5825 15484
rect 5776 15444 5782 15456
rect 5813 15453 5825 15456
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 9048 15428 9076 15524
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 6825 15419 6883 15425
rect 5644 15388 5764 15416
rect 5736 15360 5764 15388
rect 6825 15385 6837 15419
rect 6871 15416 6883 15419
rect 6914 15416 6920 15428
rect 6871 15388 6920 15416
rect 6871 15385 6883 15388
rect 6825 15379 6883 15385
rect 6914 15376 6920 15388
rect 6972 15376 6978 15428
rect 8386 15416 8392 15428
rect 8050 15388 8392 15416
rect 8386 15376 8392 15388
rect 8444 15416 8450 15428
rect 9030 15416 9036 15428
rect 8444 15388 9036 15416
rect 8444 15376 8450 15388
rect 9030 15376 9036 15388
rect 9088 15376 9094 15428
rect 9140 15416 9168 15447
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 9490 15416 9496 15428
rect 9140 15388 9496 15416
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 3234 15348 3240 15360
rect 1995 15320 3240 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 3234 15308 3240 15320
rect 3292 15348 3298 15360
rect 3970 15348 3976 15360
rect 3292 15320 3976 15348
rect 3292 15308 3298 15320
rect 3970 15308 3976 15320
rect 4028 15308 4034 15360
rect 5353 15351 5411 15357
rect 5353 15317 5365 15351
rect 5399 15348 5411 15351
rect 5718 15348 5724 15360
rect 5399 15320 5724 15348
rect 5399 15317 5411 15320
rect 5353 15311 5411 15317
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 5813 15351 5871 15357
rect 5813 15317 5825 15351
rect 5859 15348 5871 15351
rect 6454 15348 6460 15360
rect 5859 15320 6460 15348
rect 5859 15317 5871 15320
rect 5813 15311 5871 15317
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 9876 15348 9904 15524
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 11790 15552 11796 15564
rect 10275 15524 11796 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15552 12035 15555
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 12023 15524 12357 15552
rect 12023 15521 12035 15524
rect 11977 15515 12035 15521
rect 12345 15521 12357 15524
rect 12391 15552 12403 15555
rect 13081 15555 13139 15561
rect 12391 15524 13032 15552
rect 12391 15521 12403 15524
rect 12345 15515 12403 15521
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 10502 15376 10508 15428
rect 10560 15376 10566 15428
rect 10962 15416 10968 15428
rect 10888 15388 10968 15416
rect 10888 15348 10916 15388
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 12268 15416 12296 15447
rect 12710 15444 12716 15496
rect 12768 15444 12774 15496
rect 13004 15493 13032 15524
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 13127 15524 13553 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 13541 15521 13553 15524
rect 13587 15521 13599 15555
rect 16776 15552 16804 15583
rect 16776 15524 17172 15552
rect 13541 15515 13599 15521
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13446 15444 13452 15496
rect 13504 15444 13510 15496
rect 13630 15444 13636 15496
rect 13688 15444 13694 15496
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14608 15456 14657 15484
rect 14608 15444 14614 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 13648 15416 13676 15444
rect 12268 15388 13676 15416
rect 14366 15376 14372 15428
rect 14424 15416 14430 15428
rect 14844 15416 14872 15447
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 16761 15487 16819 15493
rect 16761 15484 16773 15487
rect 16172 15456 16773 15484
rect 16172 15444 16178 15456
rect 16761 15453 16773 15456
rect 16807 15453 16819 15487
rect 16761 15447 16819 15453
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 17144 15493 17172 15524
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 17310 15444 17316 15496
rect 17368 15444 17374 15496
rect 14424 15388 14872 15416
rect 14424 15376 14430 15388
rect 9876 15320 10916 15348
rect 13357 15351 13415 15357
rect 13357 15317 13369 15351
rect 13403 15348 13415 15351
rect 13814 15348 13820 15360
rect 13403 15320 13820 15348
rect 13403 15317 13415 15320
rect 13357 15311 13415 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 16945 15351 17003 15357
rect 16945 15317 16957 15351
rect 16991 15348 17003 15351
rect 17034 15348 17040 15360
rect 16991 15320 17040 15348
rect 16991 15317 17003 15320
rect 16945 15311 17003 15317
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17221 15351 17279 15357
rect 17221 15317 17233 15351
rect 17267 15348 17279 15351
rect 17586 15348 17592 15360
rect 17267 15320 17592 15348
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 1104 15258 18216 15280
rect 1104 15206 2658 15258
rect 2710 15206 2722 15258
rect 2774 15206 2786 15258
rect 2838 15206 2850 15258
rect 2902 15206 2914 15258
rect 2966 15206 2978 15258
rect 3030 15206 8658 15258
rect 8710 15206 8722 15258
rect 8774 15206 8786 15258
rect 8838 15206 8850 15258
rect 8902 15206 8914 15258
rect 8966 15206 8978 15258
rect 9030 15206 14658 15258
rect 14710 15206 14722 15258
rect 14774 15206 14786 15258
rect 14838 15206 14850 15258
rect 14902 15206 14914 15258
rect 14966 15206 14978 15258
rect 15030 15206 18216 15258
rect 1104 15184 18216 15206
rect 3970 15104 3976 15156
rect 4028 15144 4034 15156
rect 4028 15116 5488 15144
rect 4028 15104 4034 15116
rect 4062 15076 4068 15088
rect 2898 15048 4068 15076
rect 4062 15036 4068 15048
rect 4120 15076 4126 15088
rect 4120 15048 4646 15076
rect 4120 15036 4126 15048
rect 3878 14968 3884 15020
rect 3936 14968 3942 15020
rect 1394 14900 1400 14952
rect 1452 14900 1458 14952
rect 1670 14900 1676 14952
rect 1728 14900 1734 14952
rect 3896 14940 3924 14968
rect 2746 14912 3924 14940
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 2746 14804 2774 14912
rect 4154 14900 4160 14952
rect 4212 14900 4218 14952
rect 5460 14940 5488 15116
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 5592 15116 5641 15144
rect 5592 15104 5598 15116
rect 5629 15113 5641 15116
rect 5675 15113 5687 15147
rect 5629 15107 5687 15113
rect 5644 15008 5672 15107
rect 6914 15104 6920 15156
rect 6972 15104 6978 15156
rect 9306 15104 9312 15156
rect 9364 15144 9370 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9364 15116 10057 15144
rect 9364 15104 9370 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 10045 15107 10103 15113
rect 10413 15147 10471 15153
rect 10413 15113 10425 15147
rect 10459 15144 10471 15147
rect 10594 15144 10600 15156
rect 10459 15116 10600 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10594 15104 10600 15116
rect 10652 15144 10658 15156
rect 12710 15144 12716 15156
rect 10652 15116 12716 15144
rect 10652 15104 10658 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 14366 15104 14372 15156
rect 14424 15144 14430 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14424 15116 15025 15144
rect 14424 15104 14430 15116
rect 15013 15113 15025 15116
rect 15059 15144 15071 15147
rect 15657 15147 15715 15153
rect 15657 15144 15669 15147
rect 15059 15116 15669 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15657 15113 15669 15116
rect 15703 15113 15715 15147
rect 15657 15107 15715 15113
rect 9122 15036 9128 15088
rect 9180 15036 9186 15088
rect 10781 15079 10839 15085
rect 10781 15076 10793 15079
rect 10520 15048 10793 15076
rect 5905 15011 5963 15017
rect 5905 15008 5917 15011
rect 5644 14980 5917 15008
rect 5905 14977 5917 14980
rect 5951 14977 5963 15011
rect 5905 14971 5963 14977
rect 6089 15011 6147 15017
rect 6089 14977 6101 15011
rect 6135 14977 6147 15011
rect 6089 14971 6147 14977
rect 6104 14940 6132 14971
rect 6178 14968 6184 15020
rect 6236 14968 6242 15020
rect 6546 14968 6552 15020
rect 6604 14968 6610 15020
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 10520 15017 10548 15048
rect 10781 15045 10793 15048
rect 10827 15076 10839 15079
rect 11698 15076 11704 15088
rect 10827 15048 11704 15076
rect 10827 15045 10839 15048
rect 10781 15039 10839 15045
rect 11698 15036 11704 15048
rect 11756 15036 11762 15088
rect 15749 15079 15807 15085
rect 15749 15076 15761 15079
rect 15580 15048 15761 15076
rect 15580 15020 15608 15048
rect 15749 15045 15761 15048
rect 15795 15045 15807 15079
rect 15749 15039 15807 15045
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7340 14980 8217 15008
rect 7340 14968 7346 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 10229 15011 10287 15017
rect 10229 14977 10241 15011
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 14977 10655 15011
rect 10597 14971 10655 14977
rect 5460 14912 6132 14940
rect 6454 14900 6460 14952
rect 6512 14900 6518 14952
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14940 8539 14943
rect 8938 14940 8944 14952
rect 8527 14912 8944 14940
rect 8527 14909 8539 14912
rect 8481 14903 8539 14909
rect 8938 14900 8944 14912
rect 8996 14900 9002 14952
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 10244 14940 10272 14971
rect 10612 14940 10640 14971
rect 10870 14968 10876 15020
rect 10928 14968 10934 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 15008 14703 15011
rect 15102 15008 15108 15020
rect 14691 14980 15108 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 9999 14912 10640 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 10888 14872 10916 14968
rect 14550 14900 14556 14952
rect 14608 14900 14614 14952
rect 15304 14940 15332 14971
rect 15470 14968 15476 15020
rect 15528 14968 15534 15020
rect 15562 14968 15568 15020
rect 15620 14968 15626 15020
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 15930 14968 15936 15020
rect 15988 14968 15994 15020
rect 15948 14940 15976 14968
rect 15304 14912 15976 14940
rect 9732 14844 10916 14872
rect 14568 14872 14596 14900
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 14568 14844 15117 14872
rect 9732 14832 9738 14844
rect 15105 14841 15117 14844
rect 15151 14841 15163 14875
rect 15105 14835 15163 14841
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 15654 14872 15660 14884
rect 15436 14844 15660 14872
rect 15436 14832 15442 14844
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 1452 14776 2774 14804
rect 1452 14764 1458 14776
rect 3142 14764 3148 14816
rect 3200 14764 3206 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5721 14807 5779 14813
rect 5721 14804 5733 14807
rect 5684 14776 5733 14804
rect 5684 14764 5690 14776
rect 5721 14773 5733 14776
rect 5767 14773 5779 14807
rect 5721 14767 5779 14773
rect 9582 14764 9588 14816
rect 9640 14804 9646 14816
rect 10689 14807 10747 14813
rect 10689 14804 10701 14807
rect 9640 14776 10701 14804
rect 9640 14764 9646 14776
rect 10689 14773 10701 14776
rect 10735 14773 10747 14807
rect 10689 14767 10747 14773
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 1104 14714 18216 14736
rect 1104 14662 1918 14714
rect 1970 14662 1982 14714
rect 2034 14662 2046 14714
rect 2098 14662 2110 14714
rect 2162 14662 2174 14714
rect 2226 14662 2238 14714
rect 2290 14662 7918 14714
rect 7970 14662 7982 14714
rect 8034 14662 8046 14714
rect 8098 14662 8110 14714
rect 8162 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 13918 14714
rect 13970 14662 13982 14714
rect 14034 14662 14046 14714
rect 14098 14662 14110 14714
rect 14162 14662 14174 14714
rect 14226 14662 14238 14714
rect 14290 14662 18216 14714
rect 1104 14640 18216 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 1728 14572 2053 14600
rect 1728 14560 1734 14572
rect 2041 14569 2053 14572
rect 2087 14569 2099 14603
rect 2041 14563 2099 14569
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 8110 14600 8116 14612
rect 7340 14572 8116 14600
rect 7340 14560 7346 14572
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 8938 14560 8944 14612
rect 8996 14560 9002 14612
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 15930 14600 15936 14612
rect 15887 14572 15936 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 9306 14532 9312 14544
rect 9140 14504 9312 14532
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14464 2283 14467
rect 2406 14464 2412 14476
rect 2271 14436 2412 14464
rect 2271 14433 2283 14436
rect 2225 14427 2283 14433
rect 2406 14424 2412 14436
rect 2464 14464 2470 14476
rect 9140 14473 9168 14504
rect 9306 14492 9312 14504
rect 9364 14492 9370 14544
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2464 14436 2973 14464
rect 2464 14424 2470 14436
rect 2961 14433 2973 14436
rect 3007 14433 3019 14467
rect 2961 14427 3019 14433
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14433 9183 14467
rect 9125 14427 9183 14433
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 14093 14467 14151 14473
rect 14093 14433 14105 14467
rect 14139 14464 14151 14467
rect 14458 14464 14464 14476
rect 14139 14436 14464 14464
rect 14139 14433 14151 14436
rect 14093 14427 14151 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14464 17739 14467
rect 17862 14464 17868 14476
rect 17727 14436 17868 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 2314 14356 2320 14408
rect 2372 14356 2378 14408
rect 3142 14356 3148 14408
rect 3200 14356 3206 14408
rect 3418 14356 3424 14408
rect 3476 14356 3482 14408
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 4341 14399 4399 14405
rect 4341 14396 4353 14399
rect 3936 14368 4353 14396
rect 3936 14356 3942 14368
rect 4341 14365 4353 14368
rect 4387 14396 4399 14399
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4387 14368 4629 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14396 9275 14399
rect 9306 14396 9312 14408
rect 9263 14368 9312 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 6362 14288 6368 14340
rect 6420 14288 6426 14340
rect 8754 14288 8760 14340
rect 8812 14288 8818 14340
rect 11790 14288 11796 14340
rect 11848 14288 11854 14340
rect 13538 14288 13544 14340
rect 13596 14288 13602 14340
rect 14366 14288 14372 14340
rect 14424 14288 14430 14340
rect 15378 14288 15384 14340
rect 15436 14288 15442 14340
rect 15933 14331 15991 14337
rect 15933 14328 15945 14331
rect 15672 14300 15945 14328
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 2685 14263 2743 14269
rect 2685 14260 2697 14263
rect 2556 14232 2697 14260
rect 2556 14220 2562 14232
rect 2685 14229 2697 14232
rect 2731 14229 2743 14263
rect 2685 14223 2743 14229
rect 3329 14263 3387 14269
rect 3329 14229 3341 14263
rect 3375 14260 3387 14263
rect 4890 14260 4896 14272
rect 3375 14232 4896 14260
rect 3375 14229 3387 14232
rect 3329 14223 3387 14229
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 13556 14260 13584 14288
rect 15672 14260 15700 14300
rect 15933 14297 15945 14300
rect 15979 14297 15991 14331
rect 15933 14291 15991 14297
rect 13556 14232 15700 14260
rect 1104 14170 18216 14192
rect 1104 14118 2658 14170
rect 2710 14118 2722 14170
rect 2774 14118 2786 14170
rect 2838 14118 2850 14170
rect 2902 14118 2914 14170
rect 2966 14118 2978 14170
rect 3030 14118 8658 14170
rect 8710 14118 8722 14170
rect 8774 14118 8786 14170
rect 8838 14118 8850 14170
rect 8902 14118 8914 14170
rect 8966 14118 8978 14170
rect 9030 14118 14658 14170
rect 14710 14118 14722 14170
rect 14774 14118 14786 14170
rect 14838 14118 14850 14170
rect 14902 14118 14914 14170
rect 14966 14118 14978 14170
rect 15030 14118 18216 14170
rect 1104 14096 18216 14118
rect 2498 14016 2504 14068
rect 2556 14056 2562 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 2556 14028 2881 14056
rect 2556 14016 2562 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 4212 14028 5089 14056
rect 4212 14016 4218 14028
rect 5077 14025 5089 14028
rect 5123 14025 5135 14059
rect 5077 14019 5135 14025
rect 5718 14016 5724 14068
rect 5776 14016 5782 14068
rect 6365 14059 6423 14065
rect 6365 14025 6377 14059
rect 6411 14056 6423 14059
rect 6546 14056 6552 14068
rect 6411 14028 6552 14056
rect 6411 14025 6423 14028
rect 6365 14019 6423 14025
rect 2516 13988 2544 14016
rect 2516 13960 2728 13988
rect 2406 13880 2412 13932
rect 2464 13920 2470 13932
rect 2700 13929 2728 13960
rect 3142 13948 3148 14000
rect 3200 13948 3206 14000
rect 6380 13988 6408 14019
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 17770 14056 17776 14068
rect 11164 14028 11928 14056
rect 8386 13988 8392 14000
rect 5184 13960 6408 13988
rect 7406 13960 8392 13988
rect 2501 13923 2559 13929
rect 2501 13920 2513 13923
rect 2464 13892 2513 13920
rect 2464 13880 2470 13892
rect 2501 13889 2513 13892
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13889 2927 13923
rect 2869 13883 2927 13889
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3418 13920 3424 13932
rect 3007 13892 3424 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 2884 13852 2912 13883
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 4798 13852 4804 13864
rect 2884 13824 4804 13852
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5184 13852 5212 13960
rect 8386 13948 8392 13960
rect 8444 13948 8450 14000
rect 11164 13997 11192 14028
rect 11149 13991 11207 13997
rect 11149 13957 11161 13991
rect 11195 13957 11207 13991
rect 11149 13951 11207 13957
rect 11422 13948 11428 14000
rect 11480 13988 11486 14000
rect 11793 13991 11851 13997
rect 11793 13988 11805 13991
rect 11480 13960 11805 13988
rect 11480 13948 11486 13960
rect 11793 13957 11805 13960
rect 11839 13957 11851 13991
rect 11793 13951 11851 13957
rect 11900 13988 11928 14028
rect 16868 14028 17776 14056
rect 12158 13988 12164 14000
rect 11900 13960 12164 13988
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 5626 13920 5632 13932
rect 5307 13892 5632 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 8110 13880 8116 13932
rect 8168 13880 8174 13932
rect 11054 13880 11060 13932
rect 11112 13880 11118 13932
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 11296 13892 11345 13920
rect 11296 13880 11302 13892
rect 11333 13889 11345 13892
rect 11379 13889 11391 13923
rect 11333 13883 11391 13889
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 11900 13920 11928 13960
rect 12158 13948 12164 13960
rect 12216 13948 12222 14000
rect 14458 13948 14464 14000
rect 14516 13988 14522 14000
rect 16868 13997 16896 14028
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 15013 13991 15071 13997
rect 15013 13988 15025 13991
rect 14516 13960 15025 13988
rect 14516 13948 14522 13960
rect 15013 13957 15025 13960
rect 15059 13957 15071 13991
rect 15013 13951 15071 13957
rect 16853 13991 16911 13997
rect 16853 13957 16865 13991
rect 16899 13957 16911 13991
rect 16853 13951 16911 13957
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 17494 13988 17500 14000
rect 17083 13960 17500 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 17494 13948 17500 13960
rect 17552 13948 17558 14000
rect 11747 13892 11928 13920
rect 11977 13923 12035 13929
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 5184 13824 5365 13852
rect 5353 13821 5365 13824
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 7834 13812 7840 13864
rect 7892 13812 7898 13864
rect 11348 13852 11376 13883
rect 11992 13852 12020 13883
rect 11348 13824 12020 13852
rect 16776 13852 16804 13883
rect 17126 13880 17132 13932
rect 17184 13880 17190 13932
rect 17310 13880 17316 13932
rect 17368 13880 17374 13932
rect 17034 13852 17040 13864
rect 16776 13824 17040 13852
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17218 13812 17224 13864
rect 17276 13812 17282 13864
rect 2498 13676 2504 13728
rect 2556 13716 2562 13728
rect 2593 13719 2651 13725
rect 2593 13716 2605 13719
rect 2556 13688 2605 13716
rect 2556 13676 2562 13688
rect 2593 13685 2605 13688
rect 2639 13685 2651 13719
rect 2593 13679 2651 13685
rect 11241 13719 11299 13725
rect 11241 13685 11253 13719
rect 11287 13716 11299 13719
rect 11974 13716 11980 13728
rect 11287 13688 11980 13716
rect 11287 13685 11299 13688
rect 11241 13679 11299 13685
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12158 13676 12164 13728
rect 12216 13676 12222 13728
rect 16945 13719 17003 13725
rect 16945 13685 16957 13719
rect 16991 13716 17003 13719
rect 17126 13716 17132 13728
rect 16991 13688 17132 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 1104 13626 18216 13648
rect 1104 13574 1918 13626
rect 1970 13574 1982 13626
rect 2034 13574 2046 13626
rect 2098 13574 2110 13626
rect 2162 13574 2174 13626
rect 2226 13574 2238 13626
rect 2290 13574 7918 13626
rect 7970 13574 7982 13626
rect 8034 13574 8046 13626
rect 8098 13574 8110 13626
rect 8162 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 13918 13626
rect 13970 13574 13982 13626
rect 14034 13574 14046 13626
rect 14098 13574 14110 13626
rect 14162 13574 14174 13626
rect 14226 13574 14238 13626
rect 14290 13574 18216 13626
rect 1104 13552 18216 13574
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 11238 13512 11244 13524
rect 10183 13484 11244 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 11808 13484 12817 13512
rect 2498 13336 2504 13388
rect 2556 13336 2562 13388
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7282 13376 7288 13388
rect 7055 13348 7288 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13345 8815 13379
rect 8757 13339 8815 13345
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2372 13280 2421 13308
rect 2372 13268 2378 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 4798 13268 4804 13320
rect 4856 13268 4862 13320
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 4982 13308 4988 13320
rect 4939 13280 4988 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 4982 13268 4988 13280
rect 5040 13308 5046 13320
rect 5902 13308 5908 13320
rect 5040 13280 5908 13308
rect 5040 13268 5046 13280
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 8386 13268 8392 13320
rect 8444 13268 8450 13320
rect 8772 13308 8800 13339
rect 9214 13336 9220 13388
rect 9272 13336 9278 13388
rect 11808 13376 11836 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 10244 13348 11836 13376
rect 9306 13308 9312 13320
rect 8772 13280 9312 13308
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 5077 13243 5135 13249
rect 5077 13209 5089 13243
rect 5123 13240 5135 13243
rect 5350 13240 5356 13252
rect 5123 13212 5356 13240
rect 5123 13209 5135 13212
rect 5077 13203 5135 13209
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13209 7343 13243
rect 10244 13240 10272 13348
rect 12158 13336 12164 13388
rect 12216 13336 12222 13388
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12989 13379 13047 13385
rect 12989 13376 13001 13379
rect 12400 13348 13001 13376
rect 12400 13336 12406 13348
rect 12989 13345 13001 13348
rect 13035 13345 13047 13379
rect 12989 13339 13047 13345
rect 17586 13336 17592 13388
rect 17644 13336 17650 13388
rect 17862 13336 17868 13388
rect 17920 13336 17926 13388
rect 11882 13268 11888 13320
rect 11940 13268 11946 13320
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13308 12311 13311
rect 12802 13308 12808 13320
rect 12299 13280 12808 13308
rect 12299 13277 12311 13280
rect 12253 13271 12311 13277
rect 12802 13268 12808 13280
rect 12860 13308 12866 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 12860 13280 13093 13308
rect 12860 13268 12866 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 11609 13243 11667 13249
rect 7285 13203 7343 13209
rect 8864 13212 10272 13240
rect 10336 13212 10442 13240
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 2041 13175 2099 13181
rect 2041 13172 2053 13175
rect 1728 13144 2053 13172
rect 1728 13132 1734 13144
rect 2041 13141 2053 13144
rect 2087 13141 2099 13175
rect 2041 13135 2099 13141
rect 4985 13175 5043 13181
rect 4985 13141 4997 13175
rect 5031 13172 5043 13175
rect 5718 13172 5724 13184
rect 5031 13144 5724 13172
rect 5031 13141 5043 13144
rect 4985 13135 5043 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 7300 13172 7328 13203
rect 8864 13172 8892 13212
rect 7300 13144 8892 13172
rect 8941 13175 8999 13181
rect 8941 13141 8953 13175
rect 8987 13172 8999 13175
rect 9214 13172 9220 13184
rect 8987 13144 9220 13172
rect 8987 13141 8999 13144
rect 8941 13135 8999 13141
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 10336 13172 10364 13212
rect 11609 13209 11621 13243
rect 11655 13240 11667 13243
rect 11977 13243 12035 13249
rect 11977 13240 11989 13243
rect 11655 13212 11989 13240
rect 11655 13209 11667 13212
rect 11609 13203 11667 13209
rect 11977 13209 11989 13212
rect 12023 13209 12035 13243
rect 11977 13203 12035 13209
rect 15378 13200 15384 13252
rect 15436 13240 15442 13252
rect 16298 13240 16304 13252
rect 15436 13212 16304 13240
rect 15436 13200 15442 13212
rect 16298 13200 16304 13212
rect 16356 13240 16362 13252
rect 16356 13212 16422 13240
rect 16356 13200 16362 13212
rect 9640 13144 10364 13172
rect 9640 13132 9646 13144
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 12124 13144 12633 13172
rect 12124 13132 12130 13144
rect 12621 13141 12633 13144
rect 12667 13141 12679 13175
rect 12621 13135 12679 13141
rect 16117 13175 16175 13181
rect 16117 13141 16129 13175
rect 16163 13172 16175 13175
rect 16942 13172 16948 13184
rect 16163 13144 16948 13172
rect 16163 13141 16175 13144
rect 16117 13135 16175 13141
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 1104 13082 18216 13104
rect 1104 13030 2658 13082
rect 2710 13030 2722 13082
rect 2774 13030 2786 13082
rect 2838 13030 2850 13082
rect 2902 13030 2914 13082
rect 2966 13030 2978 13082
rect 3030 13030 8658 13082
rect 8710 13030 8722 13082
rect 8774 13030 8786 13082
rect 8838 13030 8850 13082
rect 8902 13030 8914 13082
rect 8966 13030 8978 13082
rect 9030 13030 14658 13082
rect 14710 13030 14722 13082
rect 14774 13030 14786 13082
rect 14838 13030 14850 13082
rect 14902 13030 14914 13082
rect 14966 13030 14978 13082
rect 15030 13030 18216 13082
rect 1104 13008 18216 13030
rect 1394 12928 1400 12980
rect 1452 12968 1458 12980
rect 1452 12940 3096 12968
rect 1452 12928 1458 12940
rect 1412 12841 1440 12928
rect 1670 12860 1676 12912
rect 1728 12860 1734 12912
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 3068 12832 3096 12940
rect 5718 12928 5724 12980
rect 5776 12928 5782 12980
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 7834 12968 7840 12980
rect 6963 12940 7840 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8444 12940 9352 12968
rect 8444 12928 8450 12940
rect 4154 12860 4160 12912
rect 4212 12860 4218 12912
rect 5534 12900 5540 12912
rect 5276 12872 5540 12900
rect 5276 12841 5304 12872
rect 5534 12860 5540 12872
rect 5592 12900 5598 12912
rect 5592 12872 6040 12900
rect 5592 12860 5598 12872
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 1397 12795 1455 12801
rect 2792 12764 2820 12818
rect 3068 12804 3249 12832
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 6012 12841 6040 12872
rect 9214 12860 9220 12912
rect 9272 12860 9278 12912
rect 9324 12900 9352 12940
rect 9582 12928 9588 12980
rect 9640 12928 9646 12980
rect 12161 12971 12219 12977
rect 12161 12937 12173 12971
rect 12207 12968 12219 12971
rect 12342 12968 12348 12980
rect 12207 12940 12348 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12802 12928 12808 12980
rect 12860 12928 12866 12980
rect 14568 12940 16436 12968
rect 9600 12900 9628 12928
rect 9324 12872 9706 12900
rect 12434 12860 12440 12912
rect 12492 12900 12498 12912
rect 12492 12872 13110 12900
rect 12492 12860 12498 12872
rect 14568 12844 14596 12940
rect 15378 12860 15384 12912
rect 15436 12860 15442 12912
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5776 12804 5825 12832
rect 5776 12792 5782 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 3513 12767 3571 12773
rect 2792 12736 3280 12764
rect 3142 12588 3148 12640
rect 3200 12588 3206 12640
rect 3252 12628 3280 12736
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 5077 12767 5135 12773
rect 5077 12764 5089 12767
rect 3559 12736 5089 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 5077 12733 5089 12736
rect 5123 12733 5135 12767
rect 5077 12727 5135 12733
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12733 5411 12767
rect 5353 12727 5411 12733
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6457 12767 6515 12773
rect 6457 12764 6469 12767
rect 5951 12736 6469 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 6457 12733 6469 12736
rect 6503 12733 6515 12767
rect 6457 12727 6515 12733
rect 5166 12656 5172 12708
rect 5224 12696 5230 12708
rect 5368 12696 5396 12727
rect 6564 12696 6592 12795
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 7340 12804 8953 12832
rect 7340 12792 7346 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 12158 12792 12164 12844
rect 12216 12792 12222 12844
rect 14550 12792 14556 12844
rect 14608 12792 14614 12844
rect 16408 12841 16436 12940
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 17405 12971 17463 12977
rect 17405 12968 17417 12971
rect 17368 12940 17417 12968
rect 17368 12928 17374 12940
rect 17405 12937 17417 12940
rect 17451 12937 17463 12971
rect 17405 12931 17463 12937
rect 16393 12835 16451 12841
rect 16393 12801 16405 12835
rect 16439 12832 16451 12835
rect 16574 12832 16580 12844
rect 16439 12804 16580 12832
rect 16439 12801 16451 12804
rect 16393 12795 16451 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12832 16911 12835
rect 17328 12832 17356 12928
rect 16899 12804 17356 12832
rect 16899 12801 16911 12804
rect 16853 12795 16911 12801
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 17552 12804 17601 12832
rect 17552 12792 17558 12804
rect 17589 12801 17601 12804
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 17770 12792 17776 12844
rect 17828 12792 17834 12844
rect 17862 12792 17868 12844
rect 17920 12792 17926 12844
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 13872 12736 14289 12764
rect 13872 12724 13878 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12764 14703 12767
rect 15102 12764 15108 12776
rect 14691 12736 15108 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 16114 12724 16120 12776
rect 16172 12724 16178 12776
rect 16942 12724 16948 12776
rect 17000 12724 17006 12776
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 17184 12736 17325 12764
rect 17184 12724 17190 12736
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 5224 12668 6592 12696
rect 5224 12656 5230 12668
rect 4154 12628 4160 12640
rect 3252 12600 4160 12628
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4985 12631 5043 12637
rect 4985 12597 4997 12631
rect 5031 12628 5043 12631
rect 5350 12628 5356 12640
rect 5031 12600 5356 12628
rect 5031 12597 5043 12600
rect 4985 12591 5043 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 10689 12631 10747 12637
rect 10689 12628 10701 12631
rect 10284 12600 10701 12628
rect 10284 12588 10290 12600
rect 10689 12597 10701 12600
rect 10735 12597 10747 12631
rect 10689 12591 10747 12597
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 1104 12538 18216 12560
rect 1104 12486 1918 12538
rect 1970 12486 1982 12538
rect 2034 12486 2046 12538
rect 2098 12486 2110 12538
rect 2162 12486 2174 12538
rect 2226 12486 2238 12538
rect 2290 12486 7918 12538
rect 7970 12486 7982 12538
rect 8034 12486 8046 12538
rect 8098 12486 8110 12538
rect 8162 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 13918 12538
rect 13970 12486 13982 12538
rect 14034 12486 14046 12538
rect 14098 12486 14110 12538
rect 14162 12486 14174 12538
rect 14226 12486 14238 12538
rect 14290 12486 18216 12538
rect 1104 12464 18216 12486
rect 5534 12384 5540 12436
rect 5592 12384 5598 12436
rect 10410 12384 10416 12436
rect 10468 12384 10474 12436
rect 16758 12424 16764 12436
rect 12406 12396 16764 12424
rect 11146 12356 11152 12368
rect 10244 12328 11152 12356
rect 4982 12180 4988 12232
rect 5040 12220 5046 12232
rect 5077 12223 5135 12229
rect 5077 12220 5089 12223
rect 5040 12192 5089 12220
rect 5040 12180 5046 12192
rect 5077 12189 5089 12192
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 5350 12180 5356 12232
rect 5408 12180 5414 12232
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7926 12220 7932 12232
rect 7156 12192 7932 12220
rect 7156 12180 7162 12192
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 8168 12192 8217 12220
rect 8168 12180 8174 12192
rect 8205 12189 8217 12192
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 8444 12192 8493 12220
rect 8444 12180 8450 12192
rect 8481 12189 8493 12192
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 8665 12223 8723 12229
rect 8665 12220 8677 12223
rect 8628 12192 8677 12220
rect 8628 12180 8634 12192
rect 8665 12189 8677 12192
rect 8711 12189 8723 12223
rect 8665 12183 8723 12189
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10244 12229 10272 12328
rect 11146 12316 11152 12328
rect 11204 12316 11210 12368
rect 11330 12288 11336 12300
rect 10612 12260 11336 12288
rect 10612 12229 10640 12260
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10192 12192 10241 12220
rect 10192 12180 10198 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 10367 12192 10609 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 10870 12180 10876 12232
rect 10928 12180 10934 12232
rect 3234 12112 3240 12164
rect 3292 12152 3298 12164
rect 6454 12152 6460 12164
rect 3292 12124 6460 12152
rect 3292 12112 3298 12124
rect 6454 12112 6460 12124
rect 6512 12152 6518 12164
rect 10505 12155 10563 12161
rect 6512 12124 10456 12152
rect 6512 12112 6518 12124
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 4614 12084 4620 12096
rect 3559 12056 4620 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 4948 12056 5181 12084
rect 4948 12044 4954 12056
rect 5169 12053 5181 12056
rect 5215 12084 5227 12087
rect 5350 12084 5356 12096
rect 5215 12056 5356 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7432 12056 8033 12084
rect 7432 12044 7438 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 10428 12084 10456 12124
rect 10505 12121 10517 12155
rect 10551 12152 10563 12155
rect 10888 12152 10916 12180
rect 12406 12152 12434 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 17494 12384 17500 12436
rect 17552 12384 17558 12436
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16574 12288 16580 12300
rect 15795 12260 16580 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 13538 12220 13544 12232
rect 12943 12192 13544 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 10551 12124 10916 12152
rect 10980 12124 12434 12152
rect 10551 12121 10563 12124
rect 10505 12115 10563 12121
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10428 12056 10701 12084
rect 10689 12053 10701 12056
rect 10735 12084 10747 12087
rect 10980 12084 11008 12124
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 13722 12152 13728 12164
rect 12768 12124 13728 12152
rect 12768 12112 12774 12124
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 16025 12155 16083 12161
rect 16025 12121 16037 12155
rect 16071 12121 16083 12155
rect 16025 12115 16083 12121
rect 10735 12056 11008 12084
rect 11057 12087 11115 12093
rect 10735 12053 10747 12056
rect 10689 12047 10747 12053
rect 11057 12053 11069 12087
rect 11103 12084 11115 12087
rect 11238 12084 11244 12096
rect 11103 12056 11244 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 13081 12087 13139 12093
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13354 12084 13360 12096
rect 13127 12056 13360 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 16040 12084 16068 12115
rect 16298 12112 16304 12164
rect 16356 12152 16362 12164
rect 16356 12124 16514 12152
rect 16356 12112 16362 12124
rect 16666 12084 16672 12096
rect 16040 12056 16672 12084
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 1104 11994 18216 12016
rect 1104 11942 2658 11994
rect 2710 11942 2722 11994
rect 2774 11942 2786 11994
rect 2838 11942 2850 11994
rect 2902 11942 2914 11994
rect 2966 11942 2978 11994
rect 3030 11942 8658 11994
rect 8710 11942 8722 11994
rect 8774 11942 8786 11994
rect 8838 11942 8850 11994
rect 8902 11942 8914 11994
rect 8966 11942 8978 11994
rect 9030 11942 14658 11994
rect 14710 11942 14722 11994
rect 14774 11942 14786 11994
rect 14838 11942 14850 11994
rect 14902 11942 14914 11994
rect 14966 11942 14978 11994
rect 15030 11942 18216 11994
rect 1104 11920 18216 11942
rect 7282 11880 7288 11892
rect 6380 11852 7288 11880
rect 1578 11772 1584 11824
rect 1636 11812 1642 11824
rect 2501 11815 2559 11821
rect 2501 11812 2513 11815
rect 1636 11784 2513 11812
rect 1636 11772 1642 11784
rect 2501 11781 2513 11784
rect 2547 11812 2559 11815
rect 2590 11812 2596 11824
rect 2547 11784 2596 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 2590 11772 2596 11784
rect 2648 11772 2654 11824
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11744 2743 11747
rect 3050 11744 3056 11756
rect 2731 11716 3056 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2424 11676 2452 11707
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3142 11704 3148 11756
rect 3200 11744 3206 11756
rect 6380 11753 6408 11852
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 8110 11840 8116 11892
rect 8168 11840 8174 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8628 11852 8861 11880
rect 8628 11840 8634 11852
rect 8849 11849 8861 11852
rect 8895 11880 8907 11883
rect 9033 11883 9091 11889
rect 9033 11880 9045 11883
rect 8895 11852 9045 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9033 11849 9045 11852
rect 9079 11849 9091 11883
rect 9033 11843 9091 11849
rect 12434 11840 12440 11892
rect 12492 11840 12498 11892
rect 13538 11840 13544 11892
rect 13596 11840 13602 11892
rect 14737 11883 14795 11889
rect 14737 11849 14749 11883
rect 14783 11880 14795 11883
rect 16114 11880 16120 11892
rect 14783 11852 16120 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 8128 11812 8156 11840
rect 8941 11815 8999 11821
rect 8941 11812 8953 11815
rect 8128 11784 8953 11812
rect 8941 11781 8953 11784
rect 8987 11781 8999 11815
rect 8941 11775 8999 11781
rect 12342 11772 12348 11824
rect 12400 11812 12406 11824
rect 12452 11812 12480 11840
rect 12400 11784 12558 11812
rect 12400 11772 12406 11784
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 3200 11716 3341 11744
rect 3200 11704 3206 11716
rect 3329 11713 3341 11716
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 8294 11744 8300 11756
rect 7774 11716 8300 11744
rect 6365 11707 6423 11713
rect 8294 11704 8300 11716
rect 8352 11704 8358 11756
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9674 11744 9680 11756
rect 9263 11716 9680 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 2372 11648 2774 11676
rect 2372 11636 2378 11648
rect 2746 11608 2774 11648
rect 3418 11636 3424 11688
rect 3476 11636 3482 11688
rect 5442 11676 5448 11688
rect 3528 11648 5448 11676
rect 3528 11608 3556 11648
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 6687 11648 8217 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8481 11679 8539 11685
rect 8481 11645 8493 11679
rect 8527 11676 8539 11679
rect 8570 11676 8576 11688
rect 8527 11648 8576 11676
rect 8527 11645 8539 11648
rect 8481 11639 8539 11645
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 2746 11580 3556 11608
rect 3694 11568 3700 11620
rect 3752 11568 3758 11620
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 9140 11608 9168 11707
rect 9674 11704 9680 11716
rect 9732 11744 9738 11756
rect 10686 11744 10692 11756
rect 9732 11716 10692 11744
rect 9732 11704 9738 11716
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 11330 11704 11336 11756
rect 11388 11704 11394 11756
rect 11790 11704 11796 11756
rect 11848 11704 11854 11756
rect 14366 11704 14372 11756
rect 14424 11704 14430 11756
rect 12066 11636 12072 11688
rect 12124 11636 12130 11688
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11676 14519 11679
rect 14734 11676 14740 11688
rect 14507 11648 14740 11676
rect 14507 11645 14519 11648
rect 14461 11639 14519 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 7984 11580 9168 11608
rect 7984 11568 7990 11580
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 10962 11608 10968 11620
rect 9640 11580 10968 11608
rect 9640 11568 9646 11580
rect 10962 11568 10968 11580
rect 11020 11568 11026 11620
rect 2593 11543 2651 11549
rect 2593 11509 2605 11543
rect 2639 11540 2651 11543
rect 2682 11540 2688 11552
rect 2639 11512 2688 11540
rect 2639 11509 2651 11512
rect 2593 11503 2651 11509
rect 2682 11500 2688 11512
rect 2740 11500 2746 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 9600 11540 9628 11568
rect 8352 11512 9628 11540
rect 8352 11500 8358 11512
rect 9858 11500 9864 11552
rect 9916 11500 9922 11552
rect 1104 11450 18216 11472
rect 1104 11398 1918 11450
rect 1970 11398 1982 11450
rect 2034 11398 2046 11450
rect 2098 11398 2110 11450
rect 2162 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 7918 11450
rect 7970 11398 7982 11450
rect 8034 11398 8046 11450
rect 8098 11398 8110 11450
rect 8162 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 13918 11450
rect 13970 11398 13982 11450
rect 14034 11398 14046 11450
rect 14098 11398 14110 11450
rect 14162 11398 14174 11450
rect 14226 11398 14238 11450
rect 14290 11398 18216 11450
rect 1104 11376 18216 11398
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5166 11336 5172 11348
rect 5031 11308 5172 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 10928 11308 11161 11336
rect 10928 11296 10934 11308
rect 11149 11305 11161 11308
rect 11195 11305 11207 11339
rect 11149 11299 11207 11305
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 12124 11308 12265 11336
rect 12124 11296 12130 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12986 11336 12992 11348
rect 12253 11299 12311 11305
rect 12820 11308 12992 11336
rect 3142 11268 3148 11280
rect 2148 11240 3148 11268
rect 2148 11132 2176 11240
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 7929 11271 7987 11277
rect 7929 11268 7941 11271
rect 6656 11240 7941 11268
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 3237 11203 3295 11209
rect 3237 11200 3249 11203
rect 2271 11172 3249 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 3237 11169 3249 11172
rect 3283 11169 3295 11203
rect 3237 11163 3295 11169
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 6656 11200 6684 11240
rect 7929 11237 7941 11240
rect 7975 11237 7987 11271
rect 7929 11231 7987 11237
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 12820 11268 12848 11308
rect 12986 11296 12992 11308
rect 13044 11336 13050 11348
rect 13044 11308 13676 11336
rect 13044 11296 13050 11308
rect 10744 11240 12848 11268
rect 10744 11228 10750 11240
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12952 11240 13185 11268
rect 12952 11228 12958 11240
rect 13173 11237 13185 11240
rect 13219 11268 13231 11271
rect 13648 11268 13676 11308
rect 14734 11296 14740 11348
rect 14792 11296 14798 11348
rect 17034 11268 17040 11280
rect 13219 11240 13584 11268
rect 13648 11240 17040 11268
rect 13219 11237 13231 11240
rect 13173 11231 13231 11237
rect 6503 11172 6684 11200
rect 6733 11203 6791 11209
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 6733 11169 6745 11203
rect 6779 11200 6791 11203
rect 7282 11200 7288 11212
rect 6779 11172 7288 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2148 11104 2329 11132
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 3050 11092 3056 11144
rect 3108 11092 3114 11144
rect 3252 11132 3280 11163
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 8478 11200 8484 11212
rect 8435 11172 8484 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 12437 11203 12495 11209
rect 10468 11172 11468 11200
rect 10468 11160 10474 11172
rect 3329 11135 3387 11141
rect 3329 11132 3341 11135
rect 3252 11104 3341 11132
rect 3329 11101 3341 11104
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11101 3571 11135
rect 3513 11095 3571 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 2700 11064 2728 11092
rect 3528 11064 3556 11095
rect 8202 11064 8208 11076
rect 2700 11036 3556 11064
rect 6026 11036 8208 11064
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 2041 10999 2099 11005
rect 2041 10996 2053 10999
rect 1728 10968 2053 10996
rect 1728 10956 1734 10968
rect 2041 10965 2053 10968
rect 2087 10965 2099 10999
rect 2041 10959 2099 10965
rect 2869 10999 2927 11005
rect 2869 10965 2881 10999
rect 2915 10996 2927 10999
rect 3142 10996 3148 11008
rect 2915 10968 3148 10996
rect 2915 10965 2927 10968
rect 2869 10959 2927 10965
rect 3142 10956 3148 10968
rect 3200 10996 3206 11008
rect 3786 10996 3792 11008
rect 3200 10968 3792 10996
rect 3200 10956 3206 10968
rect 3786 10956 3792 10968
rect 3844 10996 3850 11008
rect 4062 10996 4068 11008
rect 3844 10968 4068 10996
rect 3844 10956 3850 10968
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 6104 10996 6132 11036
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 8312 11064 8340 11095
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 9272 11104 9413 11132
rect 9272 11092 9278 11104
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 11238 11092 11244 11144
rect 11296 11092 11302 11144
rect 11440 11141 11468 11172
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 12483 11172 13400 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 13372 11144 13400 11172
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 12894 11092 12900 11144
rect 12952 11092 12958 11144
rect 12986 11092 12992 11144
rect 13044 11092 13050 11144
rect 13354 11092 13360 11144
rect 13412 11092 13418 11144
rect 13556 11141 13584 11240
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 16761 11203 16819 11209
rect 16761 11169 16773 11203
rect 16807 11200 16819 11203
rect 17218 11200 17224 11212
rect 16807 11172 17224 11200
rect 16807 11169 16819 11172
rect 16761 11163 16819 11169
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14608 11104 14657 11132
rect 14608 11092 14614 11104
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11132 14887 11135
rect 15102 11132 15108 11144
rect 14875 11104 15108 11132
rect 14875 11101 14887 11104
rect 14829 11095 14887 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 16942 11132 16948 11144
rect 16715 11104 16948 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 8478 11064 8484 11076
rect 8312 11036 8484 11064
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9674 11024 9680 11076
rect 9732 11024 9738 11076
rect 10962 11064 10968 11076
rect 10902 11036 10968 11064
rect 10962 11024 10968 11036
rect 11020 11064 11026 11076
rect 12342 11064 12348 11076
rect 11020 11036 12348 11064
rect 11020 11024 11026 11036
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 12710 11024 12716 11076
rect 12768 11064 12774 11076
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 12768 11036 13093 11064
rect 12768 11024 12774 11036
rect 13081 11033 13093 11036
rect 13127 11033 13139 11067
rect 13081 11027 13139 11033
rect 13265 11067 13323 11073
rect 13265 11033 13277 11067
rect 13311 11064 13323 11067
rect 13446 11064 13452 11076
rect 13311 11036 13452 11064
rect 13311 11033 13323 11036
rect 13265 11027 13323 11033
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 5132 10968 6132 10996
rect 5132 10956 5138 10968
rect 11238 10956 11244 11008
rect 11296 10956 11302 11008
rect 13354 10956 13360 11008
rect 13412 10956 13418 11008
rect 16301 10999 16359 11005
rect 16301 10965 16313 10999
rect 16347 10996 16359 10999
rect 16390 10996 16396 11008
rect 16347 10968 16396 10996
rect 16347 10965 16359 10968
rect 16301 10959 16359 10965
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 1104 10906 18216 10928
rect 1104 10854 2658 10906
rect 2710 10854 2722 10906
rect 2774 10854 2786 10906
rect 2838 10854 2850 10906
rect 2902 10854 2914 10906
rect 2966 10854 2978 10906
rect 3030 10854 8658 10906
rect 8710 10854 8722 10906
rect 8774 10854 8786 10906
rect 8838 10854 8850 10906
rect 8902 10854 8914 10906
rect 8966 10854 8978 10906
rect 9030 10854 14658 10906
rect 14710 10854 14722 10906
rect 14774 10854 14786 10906
rect 14838 10854 14850 10906
rect 14902 10854 14914 10906
rect 14966 10854 14978 10906
rect 15030 10854 18216 10906
rect 1104 10832 18216 10854
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3145 10795 3203 10801
rect 3145 10792 3157 10795
rect 3108 10764 3157 10792
rect 3108 10752 3114 10764
rect 3145 10761 3157 10764
rect 3191 10761 3203 10795
rect 4154 10792 4160 10804
rect 3145 10755 3203 10761
rect 3620 10764 4160 10792
rect 1670 10684 1676 10736
rect 1728 10684 1734 10736
rect 3620 10724 3648 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 9953 10795 10011 10801
rect 9953 10792 9965 10795
rect 9732 10764 9965 10792
rect 9732 10752 9738 10764
rect 9953 10761 9965 10764
rect 9999 10761 10011 10795
rect 9953 10755 10011 10761
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10468 10764 10609 10792
rect 10468 10752 10474 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 15013 10795 15071 10801
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15102 10792 15108 10804
rect 15059 10764 15108 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15102 10752 15108 10764
rect 15160 10792 15166 10804
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 15160 10764 15669 10792
rect 15160 10752 15166 10764
rect 15657 10761 15669 10764
rect 15703 10761 15715 10795
rect 15657 10755 15715 10761
rect 2898 10696 3648 10724
rect 3694 10684 3700 10736
rect 3752 10724 3758 10736
rect 4065 10727 4123 10733
rect 4065 10724 4077 10727
rect 3752 10696 4077 10724
rect 3752 10684 3758 10696
rect 4065 10693 4077 10696
rect 4111 10693 4123 10727
rect 4172 10724 4200 10752
rect 4172 10696 4554 10724
rect 4065 10687 4123 10693
rect 6454 10684 6460 10736
rect 6512 10684 6518 10736
rect 11146 10724 11152 10736
rect 10152 10696 11152 10724
rect 10152 10665 10180 10696
rect 11146 10684 11152 10696
rect 11204 10684 11210 10736
rect 15470 10724 15476 10736
rect 12406 10696 15476 10724
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10226 10616 10232 10668
rect 10284 10616 10290 10668
rect 1394 10548 1400 10600
rect 1452 10548 1458 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 2746 10560 3801 10588
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 2746 10452 2774 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 6733 10591 6791 10597
rect 6733 10588 6745 10591
rect 4120 10560 6745 10588
rect 4120 10548 4126 10560
rect 6733 10557 6745 10560
rect 6779 10588 6791 10591
rect 12406 10588 12434 10696
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 15746 10724 15752 10736
rect 15580 10696 15752 10724
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 15580 10665 15608 10696
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 17126 10724 17132 10736
rect 16546 10696 17132 10724
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14608 10628 15117 10656
rect 14608 10616 14614 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 6779 10560 12434 10588
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14424 10560 14657 10588
rect 14424 10548 14430 10560
rect 14645 10557 14657 10560
rect 14691 10588 14703 10591
rect 15304 10588 15332 10619
rect 15654 10616 15660 10668
rect 15712 10616 15718 10668
rect 15930 10616 15936 10668
rect 15988 10616 15994 10668
rect 15948 10588 15976 10616
rect 14691 10560 15148 10588
rect 15304 10560 15976 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 15120 10532 15148 10560
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 13780 10492 14596 10520
rect 13780 10480 13786 10492
rect 1452 10424 2774 10452
rect 1452 10412 1458 10424
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 5537 10455 5595 10461
rect 5537 10452 5549 10455
rect 4580 10424 5549 10452
rect 4580 10412 4586 10424
rect 5537 10421 5549 10424
rect 5583 10421 5595 10455
rect 5537 10415 5595 10421
rect 14366 10412 14372 10464
rect 14424 10412 14430 10464
rect 14568 10452 14596 10492
rect 15102 10480 15108 10532
rect 15160 10480 15166 10532
rect 16546 10452 16574 10696
rect 17126 10684 17132 10696
rect 17184 10724 17190 10736
rect 17770 10724 17776 10736
rect 17184 10696 17776 10724
rect 17184 10684 17190 10696
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 16758 10616 16764 10668
rect 16816 10616 16822 10668
rect 14568 10424 16574 10452
rect 1104 10362 18216 10384
rect 1104 10310 1918 10362
rect 1970 10310 1982 10362
rect 2034 10310 2046 10362
rect 2098 10310 2110 10362
rect 2162 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 7918 10362
rect 7970 10310 7982 10362
rect 8034 10310 8046 10362
rect 8098 10310 8110 10362
rect 8162 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 13918 10362
rect 13970 10310 13982 10362
rect 14034 10310 14046 10362
rect 14098 10310 14110 10362
rect 14162 10310 14174 10362
rect 14226 10310 14238 10362
rect 14290 10310 18216 10362
rect 1104 10288 18216 10310
rect 15654 10248 15660 10260
rect 14200 10220 15660 10248
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 6549 10183 6607 10189
rect 6549 10180 6561 10183
rect 5592 10152 6561 10180
rect 5592 10140 5598 10152
rect 6549 10149 6561 10152
rect 6595 10180 6607 10183
rect 14200 10180 14228 10220
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 15841 10251 15899 10257
rect 15841 10217 15853 10251
rect 15887 10248 15899 10251
rect 15930 10248 15936 10260
rect 15887 10220 15936 10248
rect 15887 10217 15899 10220
rect 15841 10211 15899 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 6595 10152 14228 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 5350 10112 5356 10124
rect 4724 10084 5356 10112
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 4724 10053 4752 10084
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 11238 10112 11244 10124
rect 10551 10084 11244 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 12529 10115 12587 10121
rect 12529 10081 12541 10115
rect 12575 10112 12587 10115
rect 13354 10112 13360 10124
rect 12575 10084 13360 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 14366 10072 14372 10124
rect 14424 10072 14430 10124
rect 16390 10072 16396 10124
rect 16448 10072 16454 10124
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4488 10016 4629 10044
rect 4488 10004 4494 10016
rect 4617 10013 4629 10016
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 4632 9976 4660 10007
rect 4890 10004 4896 10056
rect 4948 10004 4954 10056
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 6454 10044 6460 10056
rect 6319 10016 6460 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 6454 10004 6460 10016
rect 6512 10044 6518 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6512 10016 6837 10044
rect 6512 10004 6518 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 10226 10004 10232 10056
rect 10284 10044 10290 10056
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 10284 10016 10425 10044
rect 10284 10004 10290 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12618 10044 12624 10056
rect 12483 10016 12624 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12618 10004 12624 10016
rect 12676 10044 12682 10056
rect 13262 10044 13268 10056
rect 12676 10016 13268 10044
rect 12676 10004 12682 10016
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10013 16175 10047
rect 16117 10007 16175 10013
rect 4982 9976 4988 9988
rect 4632 9948 4988 9976
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 7193 9979 7251 9985
rect 7193 9976 7205 9979
rect 5408 9948 7205 9976
rect 5408 9936 5414 9948
rect 7193 9945 7205 9948
rect 7239 9976 7251 9979
rect 11422 9976 11428 9988
rect 7239 9948 11428 9976
rect 7239 9945 7251 9948
rect 7193 9939 7251 9945
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 5077 9911 5135 9917
rect 5077 9908 5089 9911
rect 4396 9880 5089 9908
rect 4396 9868 4402 9880
rect 5077 9877 5089 9880
rect 5123 9877 5135 9911
rect 5077 9871 5135 9877
rect 10781 9911 10839 9917
rect 10781 9877 10793 9911
rect 10827 9908 10839 9911
rect 11790 9908 11796 9920
rect 10827 9880 11796 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 12805 9911 12863 9917
rect 12805 9877 12817 9911
rect 12851 9908 12863 9911
rect 13630 9908 13636 9920
rect 12851 9880 13636 9908
rect 12851 9877 12863 9880
rect 12805 9871 12863 9877
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 14108 9908 14136 10007
rect 15378 9936 15384 9988
rect 15436 9936 15442 9988
rect 15194 9908 15200 9920
rect 14108 9880 15200 9908
rect 15194 9868 15200 9880
rect 15252 9908 15258 9920
rect 16132 9908 16160 10007
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 16540 9948 16882 9976
rect 16540 9936 16546 9948
rect 15252 9880 16160 9908
rect 15252 9868 15258 9880
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 16632 9880 17877 9908
rect 16632 9868 16638 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 1104 9818 18216 9840
rect 1104 9766 2658 9818
rect 2710 9766 2722 9818
rect 2774 9766 2786 9818
rect 2838 9766 2850 9818
rect 2902 9766 2914 9818
rect 2966 9766 2978 9818
rect 3030 9766 8658 9818
rect 8710 9766 8722 9818
rect 8774 9766 8786 9818
rect 8838 9766 8850 9818
rect 8902 9766 8914 9818
rect 8966 9766 8978 9818
rect 9030 9766 14658 9818
rect 14710 9766 14722 9818
rect 14774 9766 14786 9818
rect 14838 9766 14850 9818
rect 14902 9766 14914 9818
rect 14966 9766 14978 9818
rect 15030 9766 18216 9818
rect 1104 9744 18216 9766
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 5258 9704 5264 9716
rect 4948 9676 5264 9704
rect 4948 9664 4954 9676
rect 5258 9664 5264 9676
rect 5316 9704 5322 9716
rect 5445 9707 5503 9713
rect 5445 9704 5457 9707
rect 5316 9676 5457 9704
rect 5316 9664 5322 9676
rect 5445 9673 5457 9676
rect 5491 9673 5503 9707
rect 5445 9667 5503 9673
rect 6917 9707 6975 9713
rect 6917 9673 6929 9707
rect 6963 9673 6975 9707
rect 6917 9667 6975 9673
rect 1762 9596 1768 9648
rect 1820 9636 1826 9648
rect 2406 9636 2412 9648
rect 1820 9608 2412 9636
rect 1820 9596 1826 9608
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 6932 9636 6960 9667
rect 13262 9664 13268 9716
rect 13320 9664 13326 9716
rect 7469 9639 7527 9645
rect 7469 9636 7481 9639
rect 6932 9608 7481 9636
rect 7469 9605 7481 9608
rect 7515 9605 7527 9639
rect 7469 9599 7527 9605
rect 10045 9639 10103 9645
rect 10045 9605 10057 9639
rect 10091 9636 10103 9639
rect 10318 9636 10324 9648
rect 10091 9608 10324 9636
rect 10091 9605 10103 9608
rect 10045 9599 10103 9605
rect 10318 9596 10324 9608
rect 10376 9636 10382 9648
rect 10870 9636 10876 9648
rect 10376 9608 10876 9636
rect 10376 9596 10382 9608
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 11790 9596 11796 9648
rect 11848 9596 11854 9648
rect 12342 9596 12348 9648
rect 12400 9596 12406 9648
rect 16758 9596 16764 9648
rect 16816 9596 16822 9648
rect 17313 9639 17371 9645
rect 17313 9605 17325 9639
rect 17359 9636 17371 9639
rect 17402 9636 17408 9648
rect 17359 9608 17408 9636
rect 17359 9605 17371 9608
rect 17313 9599 17371 9605
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 2314 9528 2320 9580
rect 2372 9528 2378 9580
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 3050 9568 3056 9580
rect 2639 9540 3056 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 5074 9528 5080 9580
rect 5132 9528 5138 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 7006 9568 7012 9580
rect 6595 9540 7012 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 8570 9528 8576 9580
rect 8628 9528 8634 9580
rect 9950 9528 9956 9580
rect 10008 9528 10014 9580
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10686 9568 10692 9580
rect 10275 9540 10692 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 16776 9568 16804 9596
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 16776 9540 17233 9568
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 17494 9528 17500 9580
rect 17552 9528 17558 9580
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 3694 9500 3700 9512
rect 1452 9472 3700 9500
rect 1452 9460 1458 9472
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 3970 9460 3976 9512
rect 4028 9460 4034 9512
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 2314 9324 2320 9376
rect 2372 9324 2378 9376
rect 7208 9364 7236 9463
rect 8478 9460 8484 9512
rect 8536 9500 8542 9512
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8536 9472 8953 9500
rect 8536 9460 8542 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 9968 9500 9996 9528
rect 10134 9500 10140 9512
rect 9968 9472 10140 9500
rect 8941 9463 8999 9469
rect 10134 9460 10140 9472
rect 10192 9500 10198 9512
rect 11238 9500 11244 9512
rect 10192 9472 11244 9500
rect 10192 9460 10198 9472
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 11517 9503 11575 9509
rect 11517 9469 11529 9503
rect 11563 9500 11575 9503
rect 12434 9500 12440 9512
rect 11563 9472 12440 9500
rect 11563 9469 11575 9472
rect 11517 9463 11575 9469
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 9214 9364 9220 9376
rect 7208 9336 9220 9364
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10502 9364 10508 9376
rect 10183 9336 10508 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 17034 9324 17040 9376
rect 17092 9324 17098 9376
rect 17678 9324 17684 9376
rect 17736 9324 17742 9376
rect 1104 9274 18216 9296
rect 1104 9222 1918 9274
rect 1970 9222 1982 9274
rect 2034 9222 2046 9274
rect 2098 9222 2110 9274
rect 2162 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 7918 9274
rect 7970 9222 7982 9274
rect 8034 9222 8046 9274
rect 8098 9222 8110 9274
rect 8162 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 13918 9274
rect 13970 9222 13982 9274
rect 14034 9222 14046 9274
rect 14098 9222 14110 9274
rect 14162 9222 14174 9274
rect 14226 9222 14238 9274
rect 14290 9222 18216 9274
rect 1104 9200 18216 9222
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 6696 9132 7205 9160
rect 6696 9120 6702 9132
rect 7193 9129 7205 9132
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 8628 9132 10548 9160
rect 8628 9120 8634 9132
rect 8021 9095 8079 9101
rect 8021 9092 8033 9095
rect 7484 9064 8033 9092
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 3108 8996 3157 9024
rect 3108 8984 3114 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 5592 8996 6377 9024
rect 5592 8984 5598 8996
rect 6365 8993 6377 8996
rect 6411 8993 6423 9027
rect 6365 8987 6423 8993
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 9024 6607 9027
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 6595 8996 7389 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3752 8928 3985 8956
rect 3752 8916 3758 8928
rect 3973 8925 3985 8928
rect 4019 8956 4031 8959
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 4019 8928 4261 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 4249 8925 4261 8928
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4338 8916 4344 8968
rect 4396 8956 4402 8968
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 4396 8928 6101 8956
rect 4396 8916 4402 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 6089 8919 6147 8925
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7006 8956 7012 8968
rect 6687 8928 7012 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7116 8965 7144 8996
rect 7377 8993 7389 8996
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8956 7343 8959
rect 7484 8956 7512 9064
rect 8021 9061 8033 9064
rect 8067 9061 8079 9095
rect 8021 9055 8079 9061
rect 10520 9092 10548 9132
rect 10686 9120 10692 9172
rect 10744 9120 10750 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 15160 9132 15853 9160
rect 15160 9120 15166 9132
rect 15841 9129 15853 9132
rect 15887 9129 15899 9163
rect 15841 9123 15899 9129
rect 12342 9092 12348 9104
rect 10520 9064 12348 9092
rect 8941 9027 8999 9033
rect 7576 8996 7972 9024
rect 7576 8968 7604 8996
rect 7331 8928 7512 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 1670 8848 1676 8900
rect 1728 8848 1734 8900
rect 5074 8888 5080 8900
rect 2898 8860 5080 8888
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 5994 8848 6000 8900
rect 6052 8848 6058 8900
rect 6086 8780 6092 8832
rect 6144 8780 6150 8832
rect 7009 8823 7067 8829
rect 7009 8789 7021 8823
rect 7055 8820 7067 8823
rect 7300 8820 7328 8919
rect 7558 8916 7564 8968
rect 7616 8916 7622 8968
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7944 8965 7972 8996
rect 8941 8993 8953 9027
rect 8987 9024 8999 9027
rect 9214 9024 9220 9036
rect 8987 8996 9220 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7708 8928 7849 8956
rect 7708 8916 7714 8928
rect 7837 8925 7849 8928
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8478 8956 8484 8968
rect 8251 8928 8484 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 7852 8888 7880 8919
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 10520 8956 10548 9064
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 10928 8996 11284 9024
rect 10928 8984 10934 8996
rect 10350 8928 10548 8956
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11256 8965 11284 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 13909 9027 13967 9033
rect 13909 9024 13921 9027
rect 12492 8996 13921 9024
rect 12492 8984 12498 8996
rect 13909 8993 13921 8996
rect 13955 9024 13967 9027
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 13955 8996 14105 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 16485 9027 16543 9033
rect 16485 8993 16497 9027
rect 16531 9024 16543 9027
rect 16666 9024 16672 9036
rect 16531 8996 16672 9024
rect 16531 8993 16543 8996
rect 16485 8987 16543 8993
rect 16666 8984 16672 8996
rect 16724 9024 16730 9036
rect 17678 9024 17684 9036
rect 16724 8996 17684 9024
rect 16724 8984 16730 8996
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10744 8928 10977 8956
rect 10744 8916 10750 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 12400 8942 12558 8956
rect 12400 8928 12572 8942
rect 12400 8916 12406 8928
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 7852 8860 8125 8888
rect 8113 8857 8125 8860
rect 8159 8857 8171 8891
rect 8113 8851 8171 8857
rect 9217 8891 9275 8897
rect 9217 8857 9229 8891
rect 9263 8888 9275 8891
rect 9490 8888 9496 8900
rect 9263 8860 9496 8888
rect 9263 8857 9275 8860
rect 9217 8851 9275 8857
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 10520 8860 12204 8888
rect 7055 8792 7328 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 7745 8823 7803 8829
rect 7745 8820 7757 8823
rect 7432 8792 7757 8820
rect 7432 8780 7438 8792
rect 7745 8789 7757 8792
rect 7791 8789 7803 8823
rect 7745 8783 7803 8789
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 10520 8820 10548 8860
rect 10192 8792 10548 8820
rect 10192 8780 10198 8792
rect 10778 8780 10784 8832
rect 10836 8780 10842 8832
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 11422 8820 11428 8832
rect 11195 8792 11428 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 12176 8829 12204 8860
rect 12161 8823 12219 8829
rect 12161 8789 12173 8823
rect 12207 8789 12219 8823
rect 12544 8820 12572 8928
rect 16574 8916 16580 8968
rect 16632 8916 16638 8968
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8956 17095 8959
rect 17402 8956 17408 8968
rect 17083 8928 17408 8956
rect 17083 8925 17095 8928
rect 17037 8919 17095 8925
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 13630 8848 13636 8900
rect 13688 8848 13694 8900
rect 14366 8848 14372 8900
rect 14424 8848 14430 8900
rect 16482 8888 16488 8900
rect 14476 8860 14858 8888
rect 15672 8860 16488 8888
rect 14476 8820 14504 8860
rect 12544 8792 14504 8820
rect 14752 8820 14780 8860
rect 15378 8820 15384 8832
rect 14752 8792 15384 8820
rect 12161 8783 12219 8789
rect 15378 8780 15384 8792
rect 15436 8820 15442 8832
rect 15672 8820 15700 8860
rect 16482 8848 16488 8860
rect 16540 8888 16546 8900
rect 16758 8888 16764 8900
rect 16540 8860 16764 8888
rect 16540 8848 16546 8860
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 17126 8848 17132 8900
rect 17184 8848 17190 8900
rect 17313 8891 17371 8897
rect 17313 8857 17325 8891
rect 17359 8888 17371 8891
rect 17494 8888 17500 8900
rect 17359 8860 17500 8888
rect 17359 8857 17371 8860
rect 17313 8851 17371 8857
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 15436 8792 15700 8820
rect 15436 8780 15442 8792
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 16080 8792 16313 8820
rect 16080 8780 16086 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16301 8783 16359 8789
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 16945 8823 17003 8829
rect 16945 8820 16957 8823
rect 16908 8792 16957 8820
rect 16908 8780 16914 8792
rect 16945 8789 16957 8792
rect 16991 8820 17003 8823
rect 17037 8823 17095 8829
rect 17037 8820 17049 8823
rect 16991 8792 17049 8820
rect 16991 8789 17003 8792
rect 16945 8783 17003 8789
rect 17037 8789 17049 8792
rect 17083 8789 17095 8823
rect 17037 8783 17095 8789
rect 1104 8730 18216 8752
rect 1104 8678 2658 8730
rect 2710 8678 2722 8730
rect 2774 8678 2786 8730
rect 2838 8678 2850 8730
rect 2902 8678 2914 8730
rect 2966 8678 2978 8730
rect 3030 8678 8658 8730
rect 8710 8678 8722 8730
rect 8774 8678 8786 8730
rect 8838 8678 8850 8730
rect 8902 8678 8914 8730
rect 8966 8678 8978 8730
rect 9030 8678 14658 8730
rect 14710 8678 14722 8730
rect 14774 8678 14786 8730
rect 14838 8678 14850 8730
rect 14902 8678 14914 8730
rect 14966 8678 14978 8730
rect 15030 8678 18216 8730
rect 1104 8656 18216 8678
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3142 8616 3148 8628
rect 2915 8588 3148 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3970 8576 3976 8628
rect 4028 8616 4034 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 4028 8588 4169 8616
rect 4028 8576 4034 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 4157 8579 4215 8585
rect 4724 8588 5089 8616
rect 3050 8548 3056 8560
rect 2700 8520 3056 8548
rect 2700 8489 2728 8520
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 2976 8412 3004 8443
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 2464 8384 3004 8412
rect 4433 8415 4491 8421
rect 2464 8372 2470 8384
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4522 8412 4528 8424
rect 4479 8384 4528 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4724 8412 4752 8588
rect 5077 8585 5089 8588
rect 5123 8616 5135 8619
rect 6270 8616 6276 8628
rect 5123 8588 6276 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9548 8588 9873 8616
rect 9548 8576 9554 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 10502 8576 10508 8628
rect 10560 8576 10566 8628
rect 12621 8619 12679 8625
rect 12621 8616 12633 8619
rect 12406 8588 12633 8616
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 5258 8548 5264 8560
rect 5215 8520 5264 8548
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 5258 8508 5264 8520
rect 5316 8508 5322 8560
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4724 8384 4813 8412
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 4614 8304 4620 8356
rect 4672 8344 4678 8356
rect 4908 8344 4936 8443
rect 4982 8440 4988 8492
rect 5040 8440 5046 8492
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10520 8480 10548 8576
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 10091 8452 10456 8480
rect 10520 8452 10609 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 9950 8412 9956 8424
rect 7300 8384 9956 8412
rect 7300 8344 7328 8384
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10134 8372 10140 8424
rect 10192 8372 10198 8424
rect 10428 8412 10456 8452
rect 10597 8449 10609 8452
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 10796 8412 10824 8440
rect 10428 8384 10824 8412
rect 4672 8316 7328 8344
rect 4672 8304 4678 8316
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 9766 8344 9772 8356
rect 7432 8316 9772 8344
rect 7432 8304 7438 8316
rect 9766 8304 9772 8316
rect 9824 8344 9830 8356
rect 12406 8344 12434 8588
rect 12621 8585 12633 8588
rect 12667 8616 12679 8619
rect 13722 8616 13728 8628
rect 12667 8588 13728 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8585 15991 8619
rect 15933 8579 15991 8585
rect 15194 8548 15200 8560
rect 14476 8520 15200 8548
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 13446 8480 13452 8492
rect 12851 8452 13452 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 14476 8489 14504 8520
rect 15194 8508 15200 8520
rect 15252 8548 15258 8560
rect 15746 8548 15752 8560
rect 15252 8520 15752 8548
rect 15252 8508 15258 8520
rect 15746 8508 15752 8520
rect 15804 8548 15810 8560
rect 15948 8548 15976 8579
rect 15804 8520 15976 8548
rect 15804 8508 15810 8520
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 12544 8412 12572 8440
rect 13722 8412 13728 8424
rect 12544 8384 13728 8412
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 9824 8316 12434 8344
rect 9824 8304 9830 8316
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 17034 8344 17040 8356
rect 16724 8316 17040 8344
rect 16724 8304 16730 8316
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 2501 8279 2559 8285
rect 2501 8245 2513 8279
rect 2547 8276 2559 8279
rect 2590 8276 2596 8288
rect 2547 8248 2596 8276
rect 2547 8245 2559 8248
rect 2501 8239 2559 8245
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 10689 8279 10747 8285
rect 10689 8276 10701 8279
rect 10468 8248 10701 8276
rect 10468 8236 10474 8248
rect 10689 8245 10701 8248
rect 10735 8245 10747 8279
rect 10689 8239 10747 8245
rect 12986 8236 12992 8288
rect 13044 8236 13050 8288
rect 16761 8279 16819 8285
rect 16761 8245 16773 8279
rect 16807 8276 16819 8279
rect 16942 8276 16948 8288
rect 16807 8248 16948 8276
rect 16807 8245 16819 8248
rect 16761 8239 16819 8245
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 1104 8186 18216 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 13918 8186
rect 13970 8134 13982 8186
rect 14034 8134 14046 8186
rect 14098 8134 14110 8186
rect 14162 8134 14174 8186
rect 14226 8134 14238 8186
rect 14290 8134 18216 8186
rect 1104 8112 18216 8134
rect 1670 8032 1676 8084
rect 1728 8032 1734 8084
rect 6086 8072 6092 8084
rect 5092 8044 6092 8072
rect 2314 7896 2320 7948
rect 2372 7896 2378 7948
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 5092 7936 5120 8044
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7558 8072 7564 8084
rect 6963 8044 7564 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 12434 8032 12440 8084
rect 12492 8032 12498 8084
rect 14185 8075 14243 8081
rect 14185 8041 14197 8075
rect 14231 8072 14243 8075
rect 14366 8072 14372 8084
rect 14231 8044 14372 8072
rect 14231 8041 14243 8044
rect 14185 8035 14243 8041
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 17494 8032 17500 8084
rect 17552 8032 17558 8084
rect 4387 7908 5120 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5224 7908 7512 7936
rect 5224 7896 5230 7908
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 1872 7800 1900 7831
rect 1946 7828 1952 7880
rect 2004 7828 2010 7880
rect 2332 7868 2360 7896
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 2332 7840 2421 7868
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2590 7828 2596 7880
rect 2648 7828 2654 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4522 7868 4528 7880
rect 4295 7840 4528 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 2608 7800 2636 7828
rect 1872 7772 2636 7800
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 5534 7800 5540 7812
rect 5491 7772 5540 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 6822 7800 6828 7812
rect 6670 7772 6828 7800
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 1820 7704 2513 7732
rect 1820 7692 1826 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 4617 7735 4675 7741
rect 4617 7701 4629 7735
rect 4663 7732 4675 7735
rect 5258 7732 5264 7744
rect 4663 7704 5264 7732
rect 4663 7701 4675 7704
rect 4617 7695 4675 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 7484 7741 7512 7908
rect 14550 7896 14556 7948
rect 14608 7896 14614 7948
rect 15746 7896 15752 7948
rect 15804 7896 15810 7948
rect 16022 7896 16028 7948
rect 16080 7896 16086 7948
rect 8754 7828 8760 7880
rect 8812 7828 8818 7880
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 13909 7871 13967 7877
rect 13909 7868 13921 7871
rect 13872 7840 13921 7868
rect 13872 7828 13878 7840
rect 13909 7837 13921 7840
rect 13955 7837 13967 7871
rect 13909 7831 13967 7837
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 15764 7800 15792 7896
rect 15930 7800 15936 7812
rect 15764 7772 15936 7800
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 16758 7760 16764 7812
rect 16816 7760 16822 7812
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 9214 7732 9220 7744
rect 7515 7704 9220 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 1104 7642 18216 7664
rect 1104 7590 2658 7642
rect 2710 7590 2722 7642
rect 2774 7590 2786 7642
rect 2838 7590 2850 7642
rect 2902 7590 2914 7642
rect 2966 7590 2978 7642
rect 3030 7590 8658 7642
rect 8710 7590 8722 7642
rect 8774 7590 8786 7642
rect 8838 7590 8850 7642
rect 8902 7590 8914 7642
rect 8966 7590 8978 7642
rect 9030 7590 14658 7642
rect 14710 7590 14722 7642
rect 14774 7590 14786 7642
rect 14838 7590 14850 7642
rect 14902 7590 14914 7642
rect 14966 7590 14978 7642
rect 15030 7590 18216 7642
rect 1104 7568 18216 7590
rect 1964 7500 5580 7528
rect 1394 7284 1400 7336
rect 1452 7324 1458 7336
rect 1964 7333 1992 7500
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 4982 7460 4988 7472
rect 4856 7432 4988 7460
rect 4856 7420 4862 7432
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 5258 7420 5264 7472
rect 5316 7420 5322 7472
rect 5552 7401 5580 7500
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 6880 7500 8708 7528
rect 6880 7488 6886 7500
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 8680 7460 8708 7500
rect 9766 7488 9772 7540
rect 9824 7488 9830 7540
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14608 7500 15025 7528
rect 14608 7488 14614 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 8628 7432 8708 7460
rect 8628 7420 8634 7432
rect 9122 7420 9128 7472
rect 9180 7460 9186 7472
rect 9398 7460 9404 7472
rect 9180 7432 9404 7460
rect 9180 7420 9186 7432
rect 9398 7420 9404 7432
rect 9456 7460 9462 7472
rect 9456 7432 9904 7460
rect 9456 7420 9462 7432
rect 5537 7395 5595 7401
rect 1949 7327 2007 7333
rect 1949 7324 1961 7327
rect 1452 7296 1961 7324
rect 1452 7284 1458 7296
rect 1949 7293 1961 7296
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2314 7324 2320 7336
rect 2271 7296 2320 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 3234 7284 3240 7336
rect 3292 7324 3298 7336
rect 3344 7324 3372 7378
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 9876 7401 9904 7432
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 4798 7324 4804 7336
rect 3292 7296 4804 7324
rect 3292 7284 3298 7296
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 9600 7324 9628 7355
rect 10134 7352 10140 7404
rect 10192 7392 10198 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 10192 7364 10333 7392
rect 10192 7352 10198 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12492 7364 12541 7392
rect 12492 7352 12498 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 14737 7395 14795 7401
rect 14737 7392 14749 7395
rect 13044 7364 14749 7392
rect 13044 7352 13050 7364
rect 14737 7361 14749 7364
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 14918 7352 14924 7404
rect 14976 7352 14982 7404
rect 15010 7352 15016 7404
rect 15068 7352 15074 7404
rect 15194 7352 15200 7404
rect 15252 7352 15258 7404
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16632 7364 17049 7392
rect 16632 7352 16638 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 9324 7296 9628 7324
rect 3789 7259 3847 7265
rect 3789 7256 3801 7259
rect 3252 7228 3801 7256
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 1946 7188 1952 7200
rect 1728 7160 1952 7188
rect 1728 7148 1734 7160
rect 1946 7148 1952 7160
rect 2004 7188 2010 7200
rect 3252 7188 3280 7228
rect 3789 7225 3801 7228
rect 3835 7225 3847 7259
rect 3789 7219 3847 7225
rect 2004 7160 3280 7188
rect 2004 7148 2010 7160
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3384 7160 3709 7188
rect 3384 7148 3390 7160
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 3697 7151 3755 7157
rect 7561 7191 7619 7197
rect 7561 7157 7573 7191
rect 7607 7188 7619 7191
rect 8662 7188 8668 7200
rect 7607 7160 8668 7188
rect 7607 7157 7619 7160
rect 7561 7151 7619 7157
rect 8662 7148 8668 7160
rect 8720 7188 8726 7200
rect 9324 7188 9352 7296
rect 10410 7284 10416 7336
rect 10468 7284 10474 7336
rect 16942 7284 16948 7336
rect 17000 7284 17006 7336
rect 8720 7160 9352 7188
rect 8720 7148 8726 7160
rect 9398 7148 9404 7200
rect 9456 7148 9462 7200
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 10134 7188 10140 7200
rect 10091 7160 10140 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 14829 7191 14887 7197
rect 14829 7188 14841 7191
rect 12676 7160 14841 7188
rect 12676 7148 12682 7160
rect 14829 7157 14841 7160
rect 14875 7157 14887 7191
rect 14829 7151 14887 7157
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 1104 7098 18216 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 13918 7098
rect 13970 7046 13982 7098
rect 14034 7046 14046 7098
rect 14098 7046 14110 7098
rect 14162 7046 14174 7098
rect 14226 7046 14238 7098
rect 14290 7046 18216 7098
rect 1104 7024 18216 7046
rect 9030 6944 9036 6996
rect 9088 6984 9094 6996
rect 10134 6993 10140 6996
rect 9585 6987 9643 6993
rect 9585 6984 9597 6987
rect 9088 6956 9597 6984
rect 9088 6944 9094 6956
rect 9585 6953 9597 6956
rect 9631 6953 9643 6987
rect 9585 6947 9643 6953
rect 10124 6987 10140 6993
rect 10124 6953 10136 6987
rect 10124 6947 10140 6953
rect 10134 6944 10140 6947
rect 10192 6944 10198 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14918 6984 14924 6996
rect 13872 6956 14924 6984
rect 13872 6944 13878 6956
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15841 6987 15899 6993
rect 15841 6984 15853 6987
rect 15252 6956 15853 6984
rect 15252 6944 15258 6956
rect 15841 6953 15853 6956
rect 15887 6953 15899 6987
rect 15841 6947 15899 6953
rect 16380 6987 16438 6993
rect 16380 6953 16392 6987
rect 16426 6984 16438 6987
rect 16758 6984 16764 6996
rect 16426 6956 16764 6984
rect 16426 6953 16438 6956
rect 16380 6947 16438 6953
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 2041 6919 2099 6925
rect 2041 6885 2053 6919
rect 2087 6916 2099 6919
rect 2314 6916 2320 6928
rect 2087 6888 2320 6916
rect 2087 6885 2099 6888
rect 2041 6879 2099 6885
rect 2314 6876 2320 6888
rect 2372 6876 2378 6928
rect 15212 6916 15240 6944
rect 14936 6888 15240 6916
rect 1762 6808 1768 6860
rect 1820 6808 1826 6860
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 5224 6820 5273 6848
rect 5224 6808 5230 6820
rect 5261 6817 5273 6820
rect 5307 6817 5319 6851
rect 5261 6811 5319 6817
rect 7006 6808 7012 6860
rect 7064 6808 7070 6860
rect 9398 6848 9404 6860
rect 8404 6820 9404 6848
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 8404 6789 8432 6820
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 9907 6820 11713 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 11701 6817 11713 6820
rect 11747 6848 11759 6851
rect 12526 6848 12532 6860
rect 11747 6820 12532 6848
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 14090 6848 14096 6860
rect 13504 6820 13584 6848
rect 13504 6808 13510 6820
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 5534 6672 5540 6724
rect 5592 6672 5598 6724
rect 6822 6712 6828 6724
rect 6762 6684 6828 6712
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 8220 6712 8248 6743
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8720 6752 8769 6780
rect 8720 6740 8726 6752
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 9306 6740 9312 6792
rect 9364 6740 9370 6792
rect 13556 6789 13584 6820
rect 13648 6820 14096 6848
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 8573 6715 8631 6721
rect 8220 6684 8524 6712
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 8496 6644 8524 6684
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 9122 6712 9128 6724
rect 8619 6684 9128 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 11514 6712 11520 6724
rect 11362 6684 11520 6712
rect 11514 6672 11520 6684
rect 11572 6672 11578 6724
rect 11974 6672 11980 6724
rect 12032 6672 12038 6724
rect 13648 6712 13676 6820
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 14936 6857 14964 6888
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 14384 6820 14565 6848
rect 14384 6792 14412 6820
rect 14553 6817 14565 6820
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6848 14979 6851
rect 14967 6820 15001 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 15988 6820 16129 6848
rect 15988 6808 15994 6820
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 13202 6684 13676 6712
rect 13832 6712 13860 6743
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 15010 6780 15016 6792
rect 14507 6752 15016 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 15010 6740 15016 6752
rect 15068 6780 15074 6792
rect 15197 6783 15255 6789
rect 15197 6780 15209 6783
rect 15068 6752 15209 6780
rect 15068 6740 15074 6752
rect 15197 6749 15209 6752
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 15378 6740 15384 6792
rect 15436 6740 15442 6792
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6780 15715 6783
rect 16025 6783 16083 6789
rect 15703 6752 15884 6780
rect 15703 6749 15715 6752
rect 15657 6743 15715 6749
rect 15286 6712 15292 6724
rect 13832 6684 15292 6712
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 8496 6616 8677 6644
rect 8665 6613 8677 6616
rect 8711 6644 8723 6647
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8711 6616 8953 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 11609 6647 11667 6653
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 12250 6644 12256 6656
rect 11655 6616 12256 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 13832 6644 13860 6684
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 15396 6712 15424 6740
rect 15856 6724 15884 6752
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 16025 6743 16083 6749
rect 15749 6715 15807 6721
rect 15749 6712 15761 6715
rect 15396 6684 15761 6712
rect 15749 6681 15761 6684
rect 15795 6681 15807 6715
rect 15749 6675 15807 6681
rect 15838 6672 15844 6724
rect 15896 6712 15902 6724
rect 15933 6715 15991 6721
rect 15933 6712 15945 6715
rect 15896 6684 15945 6712
rect 15896 6672 15902 6684
rect 15933 6681 15945 6684
rect 15979 6681 15991 6715
rect 15933 6675 15991 6681
rect 16040 6712 16068 6743
rect 16482 6712 16488 6724
rect 16040 6684 16488 6712
rect 12400 6616 13860 6644
rect 12400 6604 12406 6616
rect 13998 6604 14004 6656
rect 14056 6644 14062 6656
rect 14277 6647 14335 6653
rect 14277 6644 14289 6647
rect 14056 6616 14289 6644
rect 14056 6604 14062 6616
rect 14277 6613 14289 6616
rect 14323 6613 14335 6647
rect 14277 6607 14335 6613
rect 15562 6604 15568 6656
rect 15620 6604 15626 6656
rect 15654 6604 15660 6656
rect 15712 6644 15718 6656
rect 16040 6644 16068 6684
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 16850 6672 16856 6724
rect 16908 6672 16914 6724
rect 15712 6616 16068 6644
rect 15712 6604 15718 6616
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17865 6647 17923 6653
rect 17865 6644 17877 6647
rect 17276 6616 17877 6644
rect 17276 6604 17282 6616
rect 17865 6613 17877 6616
rect 17911 6613 17923 6647
rect 17865 6607 17923 6613
rect 1104 6554 18216 6576
rect 1104 6502 2658 6554
rect 2710 6502 2722 6554
rect 2774 6502 2786 6554
rect 2838 6502 2850 6554
rect 2902 6502 2914 6554
rect 2966 6502 2978 6554
rect 3030 6502 8658 6554
rect 8710 6502 8722 6554
rect 8774 6502 8786 6554
rect 8838 6502 8850 6554
rect 8902 6502 8914 6554
rect 8966 6502 8978 6554
rect 9030 6502 14658 6554
rect 14710 6502 14722 6554
rect 14774 6502 14786 6554
rect 14838 6502 14850 6554
rect 14902 6502 14914 6554
rect 14966 6502 14978 6554
rect 15030 6502 18216 6554
rect 1104 6480 18216 6502
rect 11974 6400 11980 6452
rect 12032 6400 12038 6452
rect 12342 6440 12348 6452
rect 12084 6412 12348 6440
rect 2976 6344 3740 6372
rect 2976 6313 3004 6344
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3326 6304 3332 6316
rect 3099 6276 3332 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3712 6313 3740 6344
rect 8478 6332 8484 6384
rect 8536 6372 8542 6384
rect 12084 6372 12112 6412
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 13814 6440 13820 6452
rect 12667 6412 13820 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14148 6412 15148 6440
rect 14148 6400 14154 6412
rect 12986 6372 12992 6384
rect 8536 6344 12112 6372
rect 12406 6344 12992 6372
rect 8536 6332 8542 6344
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 3786 6304 3792 6316
rect 3743 6276 3792 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 3344 6168 3372 6264
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 3528 6236 3556 6267
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6304 12219 6307
rect 12406 6304 12434 6344
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 13998 6332 14004 6384
rect 14056 6332 14062 6384
rect 15120 6316 15148 6412
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 15473 6443 15531 6449
rect 15473 6440 15485 6443
rect 15436 6412 15485 6440
rect 15436 6400 15442 6412
rect 15473 6409 15485 6412
rect 15519 6409 15531 6443
rect 15473 6403 15531 6409
rect 15286 6332 15292 6384
rect 15344 6372 15350 6384
rect 16666 6372 16672 6384
rect 15344 6344 16672 6372
rect 15344 6332 15350 6344
rect 16666 6332 16672 6344
rect 16724 6332 16730 6384
rect 12207 6276 12434 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 12526 6264 12532 6316
rect 12584 6304 12590 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 12584 6276 13737 6304
rect 12584 6264 12590 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 16850 6304 16856 6316
rect 15160 6276 16856 6304
rect 15160 6264 15166 6276
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 3476 6208 3556 6236
rect 3476 6196 3482 6208
rect 12250 6196 12256 6248
rect 12308 6196 12314 6248
rect 15562 6236 15568 6248
rect 12406 6208 15568 6236
rect 3970 6168 3976 6180
rect 3344 6140 3976 6168
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 7558 6128 7564 6180
rect 7616 6168 7622 6180
rect 11422 6168 11428 6180
rect 7616 6140 11428 6168
rect 7616 6128 7622 6140
rect 11422 6128 11428 6140
rect 11480 6168 11486 6180
rect 12406 6168 12434 6208
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 11480 6140 12434 6168
rect 11480 6128 11486 6140
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 2777 6103 2835 6109
rect 2777 6100 2789 6103
rect 2372 6072 2789 6100
rect 2372 6060 2378 6072
rect 2777 6069 2789 6072
rect 2823 6069 2835 6103
rect 2777 6063 2835 6069
rect 3605 6103 3663 6109
rect 3605 6069 3617 6103
rect 3651 6100 3663 6103
rect 3878 6100 3884 6112
rect 3651 6072 3884 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 14090 6100 14096 6112
rect 11572 6072 14096 6100
rect 11572 6060 11578 6072
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 1104 6010 18216 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 13918 6010
rect 13970 5958 13982 6010
rect 14034 5958 14046 6010
rect 14098 5958 14110 6010
rect 14162 5958 14174 6010
rect 14226 5958 14238 6010
rect 14290 5958 18216 6010
rect 1104 5936 18216 5958
rect 3786 5856 3792 5908
rect 3844 5856 3850 5908
rect 5534 5856 5540 5908
rect 5592 5856 5598 5908
rect 7760 5868 7972 5896
rect 4614 5788 4620 5840
rect 4672 5828 4678 5840
rect 7760 5828 7788 5868
rect 4672 5800 7788 5828
rect 7837 5831 7895 5837
rect 4672 5788 4678 5800
rect 7837 5797 7849 5831
rect 7883 5797 7895 5831
rect 7837 5791 7895 5797
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1452 5732 1685 5760
rect 1452 5720 1458 5732
rect 1673 5729 1685 5732
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2314 5760 2320 5772
rect 1995 5732 2320 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 4062 5760 4068 5772
rect 3292 5732 4068 5760
rect 3292 5720 3298 5732
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5760 5411 5763
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 5399 5732 6837 5760
rect 5399 5729 5411 5732
rect 5353 5723 5411 5729
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 7006 5760 7012 5772
rect 6825 5723 6883 5729
rect 6932 5732 7012 5760
rect 1578 5652 1584 5704
rect 1636 5652 1642 5704
rect 3694 5692 3700 5704
rect 3436 5664 3700 5692
rect 3234 5624 3240 5636
rect 3174 5596 3240 5624
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 1302 5516 1308 5568
rect 1360 5556 1366 5568
rect 1397 5559 1455 5565
rect 1397 5556 1409 5559
rect 1360 5528 1409 5556
rect 1360 5516 1366 5528
rect 1397 5525 1409 5528
rect 1443 5525 1455 5559
rect 1397 5519 1455 5525
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 3326 5556 3332 5568
rect 1544 5528 3332 5556
rect 1544 5516 1550 5528
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 3436 5565 3464 5664
rect 3694 5652 3700 5664
rect 3752 5692 3758 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3752 5664 3985 5692
rect 3752 5652 3758 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 4264 5624 4292 5655
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 6932 5701 6960 5732
rect 7006 5720 7012 5732
rect 7064 5760 7070 5772
rect 7852 5760 7880 5791
rect 7064 5732 7880 5760
rect 7944 5760 7972 5868
rect 11422 5828 11428 5840
rect 10888 5800 11428 5828
rect 7944 5732 8064 5760
rect 7064 5720 7070 5732
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5661 6975 5695
rect 6917 5655 6975 5661
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 3660 5596 4292 5624
rect 3660 5584 3666 5596
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 6748 5624 6776 5655
rect 7193 5627 7251 5633
rect 7193 5624 7205 5627
rect 6604 5596 7205 5624
rect 6604 5584 6610 5596
rect 7193 5593 7205 5596
rect 7239 5593 7251 5627
rect 7392 5624 7420 5655
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 7650 5652 7656 5704
rect 7708 5692 7714 5704
rect 8036 5701 8064 5732
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 8444 5732 9229 5760
rect 8444 5720 8450 5732
rect 9217 5729 9229 5732
rect 9263 5729 9275 5763
rect 9217 5723 9275 5729
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7708 5664 7941 5692
rect 7708 5652 7714 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10652 5664 10701 5692
rect 10652 5652 10658 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 10888 5692 10916 5800
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 11146 5760 11152 5772
rect 10980 5732 11152 5760
rect 10980 5701 11008 5732
rect 11146 5720 11152 5732
rect 11204 5760 11210 5772
rect 12345 5763 12403 5769
rect 11204 5732 11560 5760
rect 11204 5720 11210 5732
rect 10827 5664 10916 5692
rect 10965 5695 11023 5701
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 10965 5661 10977 5695
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 7742 5624 7748 5636
rect 7392 5596 7748 5624
rect 7193 5587 7251 5593
rect 7742 5584 7748 5596
rect 7800 5584 7806 5636
rect 10704 5624 10732 5655
rect 11238 5652 11244 5704
rect 11296 5652 11302 5704
rect 11532 5701 11560 5732
rect 12345 5729 12357 5763
rect 12391 5760 12403 5763
rect 12618 5760 12624 5772
rect 12391 5732 12624 5760
rect 12391 5729 12403 5732
rect 12345 5723 12403 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 16025 5763 16083 5769
rect 16025 5729 16037 5763
rect 16071 5760 16083 5763
rect 17218 5760 17224 5772
rect 16071 5732 17224 5760
rect 16071 5729 16083 5732
rect 16025 5723 16083 5729
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 12250 5652 12256 5704
rect 12308 5652 12314 5704
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 16390 5692 16396 5704
rect 15979 5664 16396 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16482 5652 16488 5704
rect 16540 5652 16546 5704
rect 16574 5652 16580 5704
rect 16632 5652 16638 5704
rect 11333 5627 11391 5633
rect 11333 5624 11345 5627
rect 10704 5596 11345 5624
rect 11333 5593 11345 5596
rect 11379 5593 11391 5627
rect 11333 5587 11391 5593
rect 16758 5584 16764 5636
rect 16816 5584 16822 5636
rect 3421 5559 3479 5565
rect 3421 5525 3433 5559
rect 3467 5525 3479 5559
rect 3421 5519 3479 5525
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 7558 5556 7564 5568
rect 4203 5528 7564 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 7708 5528 8953 5556
rect 7708 5516 7714 5528
rect 8941 5525 8953 5528
rect 8987 5525 8999 5559
rect 8941 5519 8999 5525
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 11238 5556 11244 5568
rect 11195 5528 11244 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11422 5516 11428 5568
rect 11480 5516 11486 5568
rect 12621 5559 12679 5565
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 13814 5556 13820 5568
rect 12667 5528 13820 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 15102 5556 15108 5568
rect 14148 5528 15108 5556
rect 14148 5516 14154 5528
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15749 5559 15807 5565
rect 15749 5556 15761 5559
rect 15344 5528 15761 5556
rect 15344 5516 15350 5528
rect 15749 5525 15761 5528
rect 15795 5525 15807 5559
rect 15749 5519 15807 5525
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 16666 5556 16672 5568
rect 16439 5528 16672 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 1104 5466 18216 5488
rect 1104 5414 2658 5466
rect 2710 5414 2722 5466
rect 2774 5414 2786 5466
rect 2838 5414 2850 5466
rect 2902 5414 2914 5466
rect 2966 5414 2978 5466
rect 3030 5414 8658 5466
rect 8710 5414 8722 5466
rect 8774 5414 8786 5466
rect 8838 5414 8850 5466
rect 8902 5414 8914 5466
rect 8966 5414 8978 5466
rect 9030 5414 14658 5466
rect 14710 5414 14722 5466
rect 14774 5414 14786 5466
rect 14838 5414 14850 5466
rect 14902 5414 14914 5466
rect 14966 5414 14978 5466
rect 15030 5414 18216 5466
rect 1104 5392 18216 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 4614 5352 4620 5364
rect 1452 5324 3188 5352
rect 1452 5312 1458 5324
rect 2958 5284 2964 5296
rect 2438 5256 2964 5284
rect 2958 5244 2964 5256
rect 3016 5244 3022 5296
rect 3160 5225 3188 5324
rect 3252 5324 4620 5352
rect 3252 5225 3280 5324
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 7006 5312 7012 5364
rect 7064 5312 7070 5364
rect 7576 5324 9168 5352
rect 3513 5287 3571 5293
rect 3513 5253 3525 5287
rect 3559 5284 3571 5287
rect 3694 5284 3700 5296
rect 3559 5256 3700 5284
rect 3559 5253 3571 5256
rect 3513 5247 3571 5253
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 5905 5287 5963 5293
rect 4120 5256 4738 5284
rect 4120 5244 4126 5256
rect 5905 5253 5917 5287
rect 5951 5284 5963 5287
rect 7466 5284 7472 5296
rect 5951 5256 7472 5284
rect 5951 5253 5963 5256
rect 5905 5247 5963 5253
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3602 5216 3608 5228
rect 3384 5188 3608 5216
rect 3384 5176 3390 5188
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 3970 5176 3976 5228
rect 4028 5176 4034 5228
rect 7576 5225 7604 5324
rect 8294 5244 8300 5296
rect 8352 5244 8358 5296
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 6227 5188 7573 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 9140 5216 9168 5324
rect 9306 5312 9312 5364
rect 9364 5312 9370 5364
rect 11146 5312 11152 5364
rect 11204 5312 11210 5364
rect 14090 5352 14096 5364
rect 13740 5324 14096 5352
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 13740 5284 13768 5324
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 14185 5355 14243 5361
rect 14185 5321 14197 5355
rect 14231 5352 14243 5355
rect 14366 5352 14372 5364
rect 14231 5324 14372 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 16117 5355 16175 5361
rect 16117 5352 16129 5355
rect 15620 5324 16129 5352
rect 15620 5312 15626 5324
rect 16117 5321 16129 5324
rect 16163 5321 16175 5355
rect 16117 5315 16175 5321
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 16448 5324 16497 5352
rect 16448 5312 16454 5324
rect 16485 5321 16497 5324
rect 16531 5321 16543 5355
rect 16485 5315 16543 5321
rect 9272 5256 10166 5284
rect 13386 5256 13768 5284
rect 9272 5244 9278 5256
rect 13814 5244 13820 5296
rect 13872 5244 13878 5296
rect 15102 5244 15108 5296
rect 15160 5244 15166 5296
rect 16574 5284 16580 5296
rect 16040 5256 16580 5284
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9140 5188 9413 5216
rect 7561 5179 7619 5185
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1578 5148 1584 5160
rect 1443 5120 1584 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 2915 5120 3648 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3418 5040 3424 5092
rect 3476 5040 3482 5092
rect 3620 5089 3648 5120
rect 3878 5108 3884 5160
rect 3936 5108 3942 5160
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 6196 5148 6224 5179
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11020 5188 11897 5216
rect 11020 5176 11026 5188
rect 11885 5185 11897 5188
rect 11931 5216 11943 5219
rect 11931 5188 12388 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 5224 5120 6224 5148
rect 5224 5108 5230 5120
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5148 7895 5151
rect 7883 5120 9536 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 3605 5083 3663 5089
rect 3605 5049 3617 5083
rect 3651 5049 3663 5083
rect 6656 5080 6684 5111
rect 3605 5043 3663 5049
rect 6104 5052 6684 5080
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 5258 5012 5264 5024
rect 4479 4984 5264 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 5258 4972 5264 4984
rect 5316 5012 5322 5024
rect 6104 5012 6132 5052
rect 5316 4984 6132 5012
rect 5316 4972 5322 4984
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 8294 5012 8300 5024
rect 6880 4984 8300 5012
rect 6880 4972 6886 4984
rect 8294 4972 8300 4984
rect 8352 5012 8358 5024
rect 9214 5012 9220 5024
rect 8352 4984 9220 5012
rect 8352 4972 8358 4984
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9508 5012 9536 5120
rect 9674 5108 9680 5160
rect 9732 5108 9738 5160
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12360 5157 12388 5188
rect 15930 5176 15936 5228
rect 15988 5176 15994 5228
rect 16040 5225 16068 5256
rect 16574 5244 16580 5256
rect 16632 5244 16638 5296
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16758 5216 16764 5228
rect 16347 5188 16764 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 17218 5176 17224 5228
rect 17276 5176 17282 5228
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11388 5120 11805 5148
rect 11388 5108 11394 5120
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5117 12403 5151
rect 12345 5111 12403 5117
rect 14093 5151 14151 5157
rect 14093 5117 14105 5151
rect 14139 5148 14151 5151
rect 15194 5148 15200 5160
rect 14139 5120 15200 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5148 15715 5151
rect 15703 5120 16574 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 10704 5052 11529 5080
rect 10704 5012 10732 5052
rect 11517 5049 11529 5052
rect 11563 5049 11575 5083
rect 16546 5080 16574 5120
rect 17126 5108 17132 5160
rect 17184 5108 17190 5160
rect 16853 5083 16911 5089
rect 16853 5080 16865 5083
rect 16546 5052 16865 5080
rect 11517 5043 11575 5049
rect 16853 5049 16865 5052
rect 16899 5049 16911 5083
rect 16853 5043 16911 5049
rect 9508 4984 10732 5012
rect 1104 4922 18216 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 13918 4922
rect 13970 4870 13982 4922
rect 14034 4870 14046 4922
rect 14098 4870 14110 4922
rect 14162 4870 14174 4922
rect 14226 4870 14238 4922
rect 14290 4870 18216 4922
rect 1104 4848 18216 4870
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7800 4780 7849 4808
rect 7800 4768 7806 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 10505 4811 10563 4817
rect 10505 4808 10517 4811
rect 9732 4780 10517 4808
rect 9732 4768 9738 4780
rect 10505 4777 10517 4780
rect 10551 4777 10563 4811
rect 10505 4771 10563 4777
rect 11330 4768 11336 4820
rect 11388 4768 11394 4820
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 16758 4808 16764 4820
rect 16715 4780 16764 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 16853 4811 16911 4817
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 17126 4808 17132 4820
rect 16899 4780 17132 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5224 4644 6101 4672
rect 5224 4632 5230 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6362 4632 6368 4684
rect 6420 4632 6426 4684
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 11149 4675 11207 4681
rect 10735 4644 11100 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4604 10839 4607
rect 10962 4604 10968 4616
rect 10827 4576 10968 4604
rect 10827 4573 10839 4576
rect 10781 4567 10839 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11072 4604 11100 4644
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 14921 4675 14979 4681
rect 11195 4644 11468 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 11440 4616 11468 4644
rect 14921 4641 14933 4675
rect 14967 4672 14979 4675
rect 15194 4672 15200 4684
rect 14967 4644 15200 4672
rect 14967 4641 14979 4644
rect 14921 4635 14979 4641
rect 15194 4632 15200 4644
rect 15252 4672 15258 4684
rect 15930 4672 15936 4684
rect 15252 4644 15936 4672
rect 15252 4632 15258 4644
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 16448 4644 16988 4672
rect 16448 4632 16454 4644
rect 11238 4604 11244 4616
rect 11072 4576 11244 4604
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 11422 4564 11428 4616
rect 11480 4564 11486 4616
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 16960 4613 16988 4644
rect 16761 4607 16819 4613
rect 16761 4604 16773 4607
rect 16724 4576 16773 4604
rect 16724 4564 16730 4576
rect 16761 4573 16773 4576
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 6822 4496 6828 4548
rect 6880 4496 6886 4548
rect 15197 4539 15255 4545
rect 15197 4505 15209 4539
rect 15243 4536 15255 4539
rect 15286 4536 15292 4548
rect 15243 4508 15292 4536
rect 15243 4505 15255 4508
rect 15197 4499 15255 4505
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 15396 4508 15686 4536
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15396 4468 15424 4508
rect 15160 4440 15424 4468
rect 15160 4428 15166 4440
rect 1104 4378 18216 4400
rect 1104 4326 2658 4378
rect 2710 4326 2722 4378
rect 2774 4326 2786 4378
rect 2838 4326 2850 4378
rect 2902 4326 2914 4378
rect 2966 4326 2978 4378
rect 3030 4326 8658 4378
rect 8710 4326 8722 4378
rect 8774 4326 8786 4378
rect 8838 4326 8850 4378
rect 8902 4326 8914 4378
rect 8966 4326 8978 4378
rect 9030 4326 14658 4378
rect 14710 4326 14722 4378
rect 14774 4326 14786 4378
rect 14838 4326 14850 4378
rect 14902 4326 14914 4378
rect 14966 4326 14978 4378
rect 15030 4326 18216 4378
rect 1104 4304 18216 4326
rect 1104 3834 18216 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 13918 3834
rect 13970 3782 13982 3834
rect 14034 3782 14046 3834
rect 14098 3782 14110 3834
rect 14162 3782 14174 3834
rect 14226 3782 14238 3834
rect 14290 3782 18216 3834
rect 1104 3760 18216 3782
rect 1104 3290 18216 3312
rect 1104 3238 2658 3290
rect 2710 3238 2722 3290
rect 2774 3238 2786 3290
rect 2838 3238 2850 3290
rect 2902 3238 2914 3290
rect 2966 3238 2978 3290
rect 3030 3238 8658 3290
rect 8710 3238 8722 3290
rect 8774 3238 8786 3290
rect 8838 3238 8850 3290
rect 8902 3238 8914 3290
rect 8966 3238 8978 3290
rect 9030 3238 14658 3290
rect 14710 3238 14722 3290
rect 14774 3238 14786 3290
rect 14838 3238 14850 3290
rect 14902 3238 14914 3290
rect 14966 3238 14978 3290
rect 15030 3238 18216 3290
rect 1104 3216 18216 3238
rect 1104 2746 18216 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 13918 2746
rect 13970 2694 13982 2746
rect 14034 2694 14046 2746
rect 14098 2694 14110 2746
rect 14162 2694 14174 2746
rect 14226 2694 14238 2746
rect 14290 2694 18216 2746
rect 1104 2672 18216 2694
rect 15102 2456 15108 2508
rect 15160 2456 15166 2508
rect 14458 2388 14464 2440
rect 14516 2428 14522 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14516 2400 14565 2428
rect 14516 2388 14522 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 1104 2202 18216 2224
rect 1104 2150 2658 2202
rect 2710 2150 2722 2202
rect 2774 2150 2786 2202
rect 2838 2150 2850 2202
rect 2902 2150 2914 2202
rect 2966 2150 2978 2202
rect 3030 2150 8658 2202
rect 8710 2150 8722 2202
rect 8774 2150 8786 2202
rect 8838 2150 8850 2202
rect 8902 2150 8914 2202
rect 8966 2150 8978 2202
rect 9030 2150 14658 2202
rect 14710 2150 14722 2202
rect 14774 2150 14786 2202
rect 14838 2150 14850 2202
rect 14902 2150 14914 2202
rect 14966 2150 14978 2202
rect 15030 2150 18216 2202
rect 1104 2128 18216 2150
<< via1 >>
rect 1918 19014 1970 19066
rect 1982 19014 2034 19066
rect 2046 19014 2098 19066
rect 2110 19014 2162 19066
rect 2174 19014 2226 19066
rect 2238 19014 2290 19066
rect 7918 19014 7970 19066
rect 7982 19014 8034 19066
rect 8046 19014 8098 19066
rect 8110 19014 8162 19066
rect 8174 19014 8226 19066
rect 8238 19014 8290 19066
rect 13918 19014 13970 19066
rect 13982 19014 14034 19066
rect 14046 19014 14098 19066
rect 14110 19014 14162 19066
rect 14174 19014 14226 19066
rect 14238 19014 14290 19066
rect 4436 18912 4488 18964
rect 12440 18912 12492 18964
rect 1584 18844 1636 18896
rect 6828 18844 6880 18896
rect 9404 18844 9456 18896
rect 12624 18844 12676 18896
rect 1124 18708 1176 18760
rect 1676 18708 1728 18760
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 2780 18751 2832 18760
rect 2780 18717 2789 18751
rect 2789 18717 2823 18751
rect 2823 18717 2832 18751
rect 2780 18708 2832 18717
rect 5356 18776 5408 18828
rect 3148 18683 3200 18692
rect 3148 18649 3157 18683
rect 3157 18649 3191 18683
rect 3191 18649 3200 18683
rect 3148 18640 3200 18649
rect 3332 18708 3384 18760
rect 3884 18708 3936 18760
rect 4528 18751 4580 18760
rect 4528 18717 4537 18751
rect 4537 18717 4571 18751
rect 4571 18717 4580 18751
rect 4528 18708 4580 18717
rect 4988 18708 5040 18760
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 6092 18708 6144 18760
rect 6644 18708 6696 18760
rect 7288 18751 7340 18760
rect 7288 18717 7297 18751
rect 7297 18717 7331 18751
rect 7331 18717 7340 18751
rect 7288 18708 7340 18717
rect 7840 18751 7892 18760
rect 7840 18717 7849 18751
rect 7849 18717 7883 18751
rect 7883 18717 7892 18751
rect 7840 18708 7892 18717
rect 8392 18751 8444 18760
rect 8392 18717 8401 18751
rect 8401 18717 8435 18751
rect 8435 18717 8444 18751
rect 8392 18708 8444 18717
rect 8944 18751 8996 18760
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10508 18708 10560 18760
rect 11060 18708 11112 18760
rect 11612 18708 11664 18760
rect 12164 18708 12216 18760
rect 12716 18708 12768 18760
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 13820 18708 13872 18760
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 15568 18751 15620 18760
rect 15568 18717 15577 18751
rect 15577 18717 15611 18751
rect 15611 18717 15620 18751
rect 15568 18708 15620 18717
rect 16304 18751 16356 18760
rect 16304 18717 16313 18751
rect 16313 18717 16347 18751
rect 16347 18717 16356 18751
rect 16304 18708 16356 18717
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 17224 18751 17276 18760
rect 17224 18717 17233 18751
rect 17233 18717 17267 18751
rect 17267 18717 17276 18751
rect 17224 18708 17276 18717
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 1492 18572 1544 18624
rect 1768 18572 1820 18624
rect 3056 18615 3108 18624
rect 3056 18581 3065 18615
rect 3065 18581 3099 18615
rect 3099 18581 3108 18615
rect 3056 18572 3108 18581
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 3700 18572 3752 18624
rect 5172 18572 5224 18624
rect 5540 18572 5592 18624
rect 5908 18572 5960 18624
rect 7104 18572 7156 18624
rect 7472 18615 7524 18624
rect 7472 18581 7481 18615
rect 7481 18581 7515 18615
rect 7515 18581 7524 18615
rect 7472 18572 7524 18581
rect 7656 18572 7708 18624
rect 10692 18640 10744 18692
rect 10140 18572 10192 18624
rect 11336 18572 11388 18624
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 12164 18572 12216 18624
rect 12992 18615 13044 18624
rect 12992 18581 13001 18615
rect 13001 18581 13035 18615
rect 13035 18581 13044 18615
rect 12992 18572 13044 18581
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 13728 18572 13780 18624
rect 14556 18572 14608 18624
rect 15568 18572 15620 18624
rect 15752 18615 15804 18624
rect 15752 18581 15761 18615
rect 15761 18581 15795 18615
rect 15795 18581 15804 18615
rect 15752 18572 15804 18581
rect 15844 18572 15896 18624
rect 16672 18615 16724 18624
rect 16672 18581 16681 18615
rect 16681 18581 16715 18615
rect 16715 18581 16724 18615
rect 16672 18572 16724 18581
rect 17316 18572 17368 18624
rect 17776 18572 17828 18624
rect 2658 18470 2710 18522
rect 2722 18470 2774 18522
rect 2786 18470 2838 18522
rect 2850 18470 2902 18522
rect 2914 18470 2966 18522
rect 2978 18470 3030 18522
rect 8658 18470 8710 18522
rect 8722 18470 8774 18522
rect 8786 18470 8838 18522
rect 8850 18470 8902 18522
rect 8914 18470 8966 18522
rect 8978 18470 9030 18522
rect 14658 18470 14710 18522
rect 14722 18470 14774 18522
rect 14786 18470 14838 18522
rect 14850 18470 14902 18522
rect 14914 18470 14966 18522
rect 14978 18470 15030 18522
rect 3148 18411 3200 18420
rect 3148 18377 3157 18411
rect 3157 18377 3191 18411
rect 3191 18377 3200 18411
rect 3148 18368 3200 18377
rect 2412 18300 2464 18352
rect 3792 18300 3844 18352
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 2412 18164 2464 18216
rect 3148 18096 3200 18148
rect 4344 18207 4396 18216
rect 4344 18173 4353 18207
rect 4353 18173 4387 18207
rect 4387 18173 4396 18207
rect 4344 18164 4396 18173
rect 7288 18368 7340 18420
rect 8208 18368 8260 18420
rect 6920 18300 6972 18352
rect 9128 18300 9180 18352
rect 13360 18368 13412 18420
rect 13452 18368 13504 18420
rect 8208 18164 8260 18216
rect 8668 18207 8720 18216
rect 8668 18173 8677 18207
rect 8677 18173 8711 18207
rect 8711 18173 8720 18207
rect 8668 18164 8720 18173
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 13728 18343 13780 18352
rect 10600 18096 10652 18148
rect 12256 18207 12308 18216
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 13360 18275 13412 18284
rect 13360 18241 13369 18275
rect 13369 18241 13403 18275
rect 13403 18241 13412 18275
rect 13360 18232 13412 18241
rect 13728 18309 13737 18343
rect 13737 18309 13771 18343
rect 13771 18309 13780 18343
rect 13728 18300 13780 18309
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 14556 18232 14608 18284
rect 15200 18232 15252 18284
rect 15384 18164 15436 18216
rect 15936 18275 15988 18284
rect 15936 18241 15945 18275
rect 15945 18241 15979 18275
rect 15979 18241 15988 18275
rect 15936 18232 15988 18241
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 16212 18232 16264 18284
rect 18236 18232 18288 18284
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 5816 18071 5868 18080
rect 5816 18037 5825 18071
rect 5825 18037 5859 18071
rect 5859 18037 5868 18071
rect 5816 18028 5868 18037
rect 7840 18028 7892 18080
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 10416 18028 10468 18080
rect 12072 18028 12124 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 15292 18028 15344 18080
rect 16120 18096 16172 18148
rect 17592 18096 17644 18148
rect 15660 18071 15712 18080
rect 15660 18037 15669 18071
rect 15669 18037 15703 18071
rect 15703 18037 15712 18071
rect 15660 18028 15712 18037
rect 15936 18028 15988 18080
rect 17684 18071 17736 18080
rect 17684 18037 17693 18071
rect 17693 18037 17727 18071
rect 17727 18037 17736 18071
rect 17684 18028 17736 18037
rect 1918 17926 1970 17978
rect 1982 17926 2034 17978
rect 2046 17926 2098 17978
rect 2110 17926 2162 17978
rect 2174 17926 2226 17978
rect 2238 17926 2290 17978
rect 7918 17926 7970 17978
rect 7982 17926 8034 17978
rect 8046 17926 8098 17978
rect 8110 17926 8162 17978
rect 8174 17926 8226 17978
rect 8238 17926 8290 17978
rect 13918 17926 13970 17978
rect 13982 17926 14034 17978
rect 14046 17926 14098 17978
rect 14110 17926 14162 17978
rect 14174 17926 14226 17978
rect 14238 17926 14290 17978
rect 1676 17824 1728 17876
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 8668 17824 8720 17876
rect 5264 17756 5316 17808
rect 2504 17688 2556 17740
rect 3056 17731 3108 17740
rect 3056 17697 3065 17731
rect 3065 17697 3099 17731
rect 3099 17697 3108 17731
rect 3056 17688 3108 17697
rect 3240 17620 3292 17672
rect 5172 17620 5224 17672
rect 3792 17552 3844 17604
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 7748 17688 7800 17740
rect 12808 17824 12860 17876
rect 13544 17867 13596 17876
rect 13544 17833 13553 17867
rect 13553 17833 13587 17867
rect 13587 17833 13596 17867
rect 13544 17824 13596 17833
rect 15200 17824 15252 17876
rect 12072 17731 12124 17740
rect 12072 17697 12081 17731
rect 12081 17697 12115 17731
rect 12115 17697 12124 17731
rect 12072 17688 12124 17697
rect 14556 17688 14608 17740
rect 17868 17731 17920 17740
rect 17868 17697 17877 17731
rect 17877 17697 17911 17731
rect 17911 17697 17920 17731
rect 17868 17688 17920 17697
rect 5816 17620 5868 17672
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 4620 17484 4672 17536
rect 6828 17552 6880 17604
rect 7840 17620 7892 17672
rect 9772 17663 9824 17672
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 10416 17663 10468 17672
rect 10416 17629 10425 17663
rect 10425 17629 10459 17663
rect 10459 17629 10468 17663
rect 10416 17620 10468 17629
rect 11612 17620 11664 17672
rect 13820 17552 13872 17604
rect 15476 17552 15528 17604
rect 16304 17552 16356 17604
rect 17592 17595 17644 17604
rect 17592 17561 17601 17595
rect 17601 17561 17635 17595
rect 17635 17561 17644 17595
rect 17592 17552 17644 17561
rect 10232 17527 10284 17536
rect 10232 17493 10241 17527
rect 10241 17493 10275 17527
rect 10275 17493 10284 17527
rect 10232 17484 10284 17493
rect 11152 17527 11204 17536
rect 11152 17493 11161 17527
rect 11161 17493 11195 17527
rect 11195 17493 11204 17527
rect 11152 17484 11204 17493
rect 12256 17484 12308 17536
rect 2658 17382 2710 17434
rect 2722 17382 2774 17434
rect 2786 17382 2838 17434
rect 2850 17382 2902 17434
rect 2914 17382 2966 17434
rect 2978 17382 3030 17434
rect 8658 17382 8710 17434
rect 8722 17382 8774 17434
rect 8786 17382 8838 17434
rect 8850 17382 8902 17434
rect 8914 17382 8966 17434
rect 8978 17382 9030 17434
rect 14658 17382 14710 17434
rect 14722 17382 14774 17434
rect 14786 17382 14838 17434
rect 14850 17382 14902 17434
rect 14914 17382 14966 17434
rect 14978 17382 15030 17434
rect 4344 17280 4396 17332
rect 7564 17280 7616 17332
rect 9772 17280 9824 17332
rect 15476 17323 15528 17332
rect 15476 17289 15485 17323
rect 15485 17289 15519 17323
rect 15519 17289 15528 17323
rect 15476 17280 15528 17289
rect 6828 17212 6880 17264
rect 1400 17144 1452 17196
rect 2504 17144 2556 17196
rect 4620 17187 4672 17196
rect 4620 17153 4629 17187
rect 4629 17153 4663 17187
rect 4663 17153 4672 17187
rect 4620 17144 4672 17153
rect 5264 17144 5316 17196
rect 7748 17212 7800 17264
rect 9128 17212 9180 17264
rect 11152 17212 11204 17264
rect 15660 17212 15712 17264
rect 3240 17076 3292 17128
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 4252 17008 4304 17060
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 7748 17076 7800 17128
rect 11520 17076 11572 17128
rect 16212 17076 16264 17128
rect 4804 16940 4856 16992
rect 7656 16940 7708 16992
rect 10876 16940 10928 16992
rect 1918 16838 1970 16890
rect 1982 16838 2034 16890
rect 2046 16838 2098 16890
rect 2110 16838 2162 16890
rect 2174 16838 2226 16890
rect 2238 16838 2290 16890
rect 7918 16838 7970 16890
rect 7982 16838 8034 16890
rect 8046 16838 8098 16890
rect 8110 16838 8162 16890
rect 8174 16838 8226 16890
rect 8238 16838 8290 16890
rect 13918 16838 13970 16890
rect 13982 16838 14034 16890
rect 14046 16838 14098 16890
rect 14110 16838 14162 16890
rect 14174 16838 14226 16890
rect 14238 16838 14290 16890
rect 1400 16779 1452 16788
rect 1400 16745 1409 16779
rect 1409 16745 1443 16779
rect 1443 16745 1452 16779
rect 1400 16736 1452 16745
rect 16212 16736 16264 16788
rect 3148 16643 3200 16652
rect 3148 16609 3157 16643
rect 3157 16609 3191 16643
rect 3191 16609 3200 16643
rect 3148 16600 3200 16609
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 7288 16600 7340 16652
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 10232 16600 10284 16652
rect 10876 16600 10928 16652
rect 4712 16532 4764 16541
rect 7196 16532 7248 16584
rect 7840 16532 7892 16584
rect 9772 16532 9824 16584
rect 14556 16600 14608 16652
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 13084 16532 13136 16584
rect 2412 16464 2464 16516
rect 4068 16464 4120 16516
rect 13268 16464 13320 16516
rect 14188 16464 14240 16516
rect 10508 16396 10560 16448
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 13820 16396 13872 16448
rect 15292 16396 15344 16448
rect 16304 16464 16356 16516
rect 17592 16507 17644 16516
rect 17592 16473 17601 16507
rect 17601 16473 17635 16507
rect 17635 16473 17644 16507
rect 17592 16464 17644 16473
rect 16120 16439 16172 16448
rect 16120 16405 16129 16439
rect 16129 16405 16163 16439
rect 16163 16405 16172 16439
rect 16120 16396 16172 16405
rect 2658 16294 2710 16346
rect 2722 16294 2774 16346
rect 2786 16294 2838 16346
rect 2850 16294 2902 16346
rect 2914 16294 2966 16346
rect 2978 16294 3030 16346
rect 8658 16294 8710 16346
rect 8722 16294 8774 16346
rect 8786 16294 8838 16346
rect 8850 16294 8902 16346
rect 8914 16294 8966 16346
rect 8978 16294 9030 16346
rect 14658 16294 14710 16346
rect 14722 16294 14774 16346
rect 14786 16294 14838 16346
rect 14850 16294 14902 16346
rect 14914 16294 14966 16346
rect 14978 16294 15030 16346
rect 4068 16192 4120 16244
rect 4252 16167 4304 16176
rect 4252 16133 4261 16167
rect 4261 16133 4295 16167
rect 4295 16133 4304 16167
rect 4252 16124 4304 16133
rect 11060 16124 11112 16176
rect 13820 16192 13872 16244
rect 14188 16235 14240 16244
rect 14188 16201 14197 16235
rect 14197 16201 14231 16235
rect 14231 16201 14240 16235
rect 14188 16192 14240 16201
rect 16120 16192 16172 16244
rect 13268 16124 13320 16176
rect 3240 15988 3292 16040
rect 3884 15988 3936 16040
rect 13084 16056 13136 16108
rect 13452 16099 13504 16108
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 16764 16124 16816 16176
rect 13452 16056 13504 16065
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 2320 15852 2372 15904
rect 11888 15988 11940 16040
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 15108 16056 15160 16108
rect 14740 15988 14792 16040
rect 15476 15920 15528 15972
rect 17684 16124 17736 16176
rect 11796 15852 11848 15904
rect 13636 15852 13688 15904
rect 17040 15852 17092 15904
rect 17316 15852 17368 15904
rect 17592 15852 17644 15904
rect 1918 15750 1970 15802
rect 1982 15750 2034 15802
rect 2046 15750 2098 15802
rect 2110 15750 2162 15802
rect 2174 15750 2226 15802
rect 2238 15750 2290 15802
rect 7918 15750 7970 15802
rect 7982 15750 8034 15802
rect 8046 15750 8098 15802
rect 8110 15750 8162 15802
rect 8174 15750 8226 15802
rect 8238 15750 8290 15802
rect 13918 15750 13970 15802
rect 13982 15750 14034 15802
rect 14046 15750 14098 15802
rect 14110 15750 14162 15802
rect 14174 15750 14226 15802
rect 14238 15750 14290 15802
rect 7840 15648 7892 15700
rect 11888 15648 11940 15700
rect 14740 15691 14792 15700
rect 14740 15657 14749 15691
rect 14749 15657 14783 15691
rect 14783 15657 14792 15691
rect 14740 15648 14792 15657
rect 12716 15580 12768 15632
rect 13452 15580 13504 15632
rect 5540 15512 5592 15564
rect 6184 15512 6236 15564
rect 7288 15512 7340 15564
rect 940 15444 992 15496
rect 4804 15444 4856 15496
rect 5540 15376 5592 15428
rect 5724 15444 5776 15496
rect 6920 15376 6972 15428
rect 8392 15376 8444 15428
rect 9036 15376 9088 15428
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 9496 15376 9548 15428
rect 3240 15308 3292 15360
rect 3976 15308 4028 15360
rect 5724 15308 5776 15360
rect 6460 15308 6512 15360
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 11796 15512 11848 15564
rect 10508 15419 10560 15428
rect 10508 15385 10517 15419
rect 10517 15385 10551 15419
rect 10551 15385 10560 15419
rect 10508 15376 10560 15385
rect 10968 15376 11020 15428
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 14556 15444 14608 15496
rect 14372 15376 14424 15428
rect 16120 15444 16172 15496
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 13820 15308 13872 15360
rect 17040 15308 17092 15360
rect 17592 15308 17644 15360
rect 2658 15206 2710 15258
rect 2722 15206 2774 15258
rect 2786 15206 2838 15258
rect 2850 15206 2902 15258
rect 2914 15206 2966 15258
rect 2978 15206 3030 15258
rect 8658 15206 8710 15258
rect 8722 15206 8774 15258
rect 8786 15206 8838 15258
rect 8850 15206 8902 15258
rect 8914 15206 8966 15258
rect 8978 15206 9030 15258
rect 14658 15206 14710 15258
rect 14722 15206 14774 15258
rect 14786 15206 14838 15258
rect 14850 15206 14902 15258
rect 14914 15206 14966 15258
rect 14978 15206 15030 15258
rect 3976 15104 4028 15156
rect 4068 15036 4120 15088
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 1400 14764 1452 14816
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 5540 15104 5592 15156
rect 6920 15147 6972 15156
rect 6920 15113 6929 15147
rect 6929 15113 6963 15147
rect 6963 15113 6972 15147
rect 6920 15104 6972 15113
rect 9312 15104 9364 15156
rect 10600 15104 10652 15156
rect 12716 15104 12768 15156
rect 14372 15104 14424 15156
rect 9128 15036 9180 15088
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 7288 14968 7340 15020
rect 11704 15036 11756 15088
rect 6460 14943 6512 14952
rect 6460 14909 6469 14943
rect 6469 14909 6503 14943
rect 6503 14909 6512 14943
rect 6460 14900 6512 14909
rect 8944 14900 8996 14952
rect 10876 15011 10928 15020
rect 10876 14977 10885 15011
rect 10885 14977 10919 15011
rect 10919 14977 10928 15011
rect 10876 14968 10928 14977
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 15108 14968 15160 15020
rect 9680 14832 9732 14884
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 15936 15011 15988 15020
rect 15936 14977 15945 15011
rect 15945 14977 15979 15011
rect 15979 14977 15988 15011
rect 15936 14968 15988 14977
rect 15384 14832 15436 14884
rect 15660 14832 15712 14884
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 5632 14764 5684 14816
rect 9588 14764 9640 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 1918 14662 1970 14714
rect 1982 14662 2034 14714
rect 2046 14662 2098 14714
rect 2110 14662 2162 14714
rect 2174 14662 2226 14714
rect 2238 14662 2290 14714
rect 7918 14662 7970 14714
rect 7982 14662 8034 14714
rect 8046 14662 8098 14714
rect 8110 14662 8162 14714
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 13918 14662 13970 14714
rect 13982 14662 14034 14714
rect 14046 14662 14098 14714
rect 14110 14662 14162 14714
rect 14174 14662 14226 14714
rect 14238 14662 14290 14714
rect 1676 14560 1728 14612
rect 7288 14603 7340 14612
rect 7288 14569 7297 14603
rect 7297 14569 7331 14603
rect 7331 14569 7340 14603
rect 7288 14560 7340 14569
rect 8116 14560 8168 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 15936 14560 15988 14612
rect 2412 14424 2464 14476
rect 9312 14492 9364 14544
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 14464 14424 14516 14476
rect 17868 14424 17920 14476
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 3884 14356 3936 14408
rect 9312 14356 9364 14408
rect 6368 14331 6420 14340
rect 6368 14297 6377 14331
rect 6377 14297 6411 14331
rect 6411 14297 6420 14331
rect 6368 14288 6420 14297
rect 8760 14331 8812 14340
rect 8760 14297 8769 14331
rect 8769 14297 8803 14331
rect 8803 14297 8812 14331
rect 8760 14288 8812 14297
rect 11796 14331 11848 14340
rect 11796 14297 11805 14331
rect 11805 14297 11839 14331
rect 11839 14297 11848 14331
rect 11796 14288 11848 14297
rect 13544 14331 13596 14340
rect 13544 14297 13553 14331
rect 13553 14297 13587 14331
rect 13587 14297 13596 14331
rect 13544 14288 13596 14297
rect 14372 14331 14424 14340
rect 14372 14297 14381 14331
rect 14381 14297 14415 14331
rect 14415 14297 14424 14331
rect 14372 14288 14424 14297
rect 15384 14288 15436 14340
rect 2504 14220 2556 14272
rect 4896 14220 4948 14272
rect 2658 14118 2710 14170
rect 2722 14118 2774 14170
rect 2786 14118 2838 14170
rect 2850 14118 2902 14170
rect 2914 14118 2966 14170
rect 2978 14118 3030 14170
rect 8658 14118 8710 14170
rect 8722 14118 8774 14170
rect 8786 14118 8838 14170
rect 8850 14118 8902 14170
rect 8914 14118 8966 14170
rect 8978 14118 9030 14170
rect 14658 14118 14710 14170
rect 14722 14118 14774 14170
rect 14786 14118 14838 14170
rect 14850 14118 14902 14170
rect 14914 14118 14966 14170
rect 14978 14118 15030 14170
rect 2504 14016 2556 14068
rect 4160 14016 4212 14068
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 2412 13880 2464 13932
rect 3148 13991 3200 14000
rect 3148 13957 3157 13991
rect 3157 13957 3191 13991
rect 3191 13957 3200 13991
rect 3148 13948 3200 13957
rect 6552 14016 6604 14068
rect 3424 13880 3476 13932
rect 4804 13812 4856 13864
rect 8392 13948 8444 14000
rect 11428 13948 11480 14000
rect 5632 13880 5684 13932
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 11244 13880 11296 13932
rect 12164 13948 12216 14000
rect 14464 13948 14516 14000
rect 17776 14016 17828 14068
rect 17500 13948 17552 14000
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 17316 13923 17368 13932
rect 17316 13889 17325 13923
rect 17325 13889 17359 13923
rect 17359 13889 17368 13923
rect 17316 13880 17368 13889
rect 17040 13812 17092 13864
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 2504 13676 2556 13728
rect 11980 13676 12032 13728
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 12164 13676 12216 13685
rect 17132 13676 17184 13728
rect 1918 13574 1970 13626
rect 1982 13574 2034 13626
rect 2046 13574 2098 13626
rect 2110 13574 2162 13626
rect 2174 13574 2226 13626
rect 2238 13574 2290 13626
rect 7918 13574 7970 13626
rect 7982 13574 8034 13626
rect 8046 13574 8098 13626
rect 8110 13574 8162 13626
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 13918 13574 13970 13626
rect 13982 13574 14034 13626
rect 14046 13574 14098 13626
rect 14110 13574 14162 13626
rect 14174 13574 14226 13626
rect 14238 13574 14290 13626
rect 11244 13472 11296 13524
rect 2504 13379 2556 13388
rect 2504 13345 2513 13379
rect 2513 13345 2547 13379
rect 2547 13345 2556 13379
rect 2504 13336 2556 13345
rect 7288 13336 7340 13388
rect 2320 13268 2372 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 4988 13268 5040 13320
rect 5908 13268 5960 13320
rect 8392 13268 8444 13320
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 5356 13200 5408 13252
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 12348 13336 12400 13388
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 17868 13379 17920 13388
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 11888 13311 11940 13320
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 12808 13268 12860 13320
rect 1676 13132 1728 13184
rect 5724 13132 5776 13184
rect 9220 13132 9272 13184
rect 9588 13132 9640 13184
rect 15384 13200 15436 13252
rect 16304 13200 16356 13252
rect 12072 13132 12124 13184
rect 16948 13132 17000 13184
rect 2658 13030 2710 13082
rect 2722 13030 2774 13082
rect 2786 13030 2838 13082
rect 2850 13030 2902 13082
rect 2914 13030 2966 13082
rect 2978 13030 3030 13082
rect 8658 13030 8710 13082
rect 8722 13030 8774 13082
rect 8786 13030 8838 13082
rect 8850 13030 8902 13082
rect 8914 13030 8966 13082
rect 8978 13030 9030 13082
rect 14658 13030 14710 13082
rect 14722 13030 14774 13082
rect 14786 13030 14838 13082
rect 14850 13030 14902 13082
rect 14914 13030 14966 13082
rect 14978 13030 15030 13082
rect 1400 12928 1452 12980
rect 1676 12903 1728 12912
rect 1676 12869 1685 12903
rect 1685 12869 1719 12903
rect 1719 12869 1728 12903
rect 1676 12860 1728 12869
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 7840 12928 7892 12980
rect 8392 12928 8444 12980
rect 4160 12860 4212 12912
rect 5540 12860 5592 12912
rect 5724 12792 5776 12844
rect 9220 12903 9272 12912
rect 9220 12869 9229 12903
rect 9229 12869 9263 12903
rect 9263 12869 9272 12903
rect 9220 12860 9272 12869
rect 9588 12928 9640 12980
rect 12348 12928 12400 12980
rect 12808 12971 12860 12980
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 12440 12860 12492 12912
rect 15384 12860 15436 12912
rect 3148 12631 3200 12640
rect 3148 12597 3157 12631
rect 3157 12597 3191 12631
rect 3191 12597 3200 12631
rect 3148 12588 3200 12597
rect 5172 12656 5224 12708
rect 7288 12792 7340 12844
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 12164 12835 12216 12844
rect 12164 12801 12173 12835
rect 12173 12801 12207 12835
rect 12207 12801 12216 12835
rect 12164 12792 12216 12801
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 17316 12928 17368 12980
rect 16580 12792 16632 12844
rect 17500 12792 17552 12844
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 13820 12724 13872 12776
rect 15108 12724 15160 12776
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 16120 12724 16172 12733
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 17132 12724 17184 12776
rect 4160 12588 4212 12640
rect 5356 12588 5408 12640
rect 10232 12588 10284 12640
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 1918 12486 1970 12538
rect 1982 12486 2034 12538
rect 2046 12486 2098 12538
rect 2110 12486 2162 12538
rect 2174 12486 2226 12538
rect 2238 12486 2290 12538
rect 7918 12486 7970 12538
rect 7982 12486 8034 12538
rect 8046 12486 8098 12538
rect 8110 12486 8162 12538
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 13918 12486 13970 12538
rect 13982 12486 14034 12538
rect 14046 12486 14098 12538
rect 14110 12486 14162 12538
rect 14174 12486 14226 12538
rect 14238 12486 14290 12538
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 10416 12427 10468 12436
rect 10416 12393 10425 12427
rect 10425 12393 10459 12427
rect 10459 12393 10468 12427
rect 10416 12384 10468 12393
rect 4988 12180 5040 12232
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 7104 12180 7156 12232
rect 7932 12223 7984 12232
rect 7932 12189 7941 12223
rect 7941 12189 7975 12223
rect 7975 12189 7984 12223
rect 7932 12180 7984 12189
rect 8116 12180 8168 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8576 12180 8628 12232
rect 10140 12180 10192 12232
rect 11152 12316 11204 12368
rect 11336 12248 11388 12300
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 3240 12155 3292 12164
rect 3240 12121 3249 12155
rect 3249 12121 3283 12155
rect 3283 12121 3292 12155
rect 3240 12112 3292 12121
rect 6460 12112 6512 12164
rect 4620 12044 4672 12096
rect 4896 12044 4948 12096
rect 5356 12044 5408 12096
rect 7380 12044 7432 12096
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 16764 12384 16816 12436
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 16580 12248 16632 12300
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 13544 12180 13596 12232
rect 12716 12155 12768 12164
rect 12716 12121 12725 12155
rect 12725 12121 12759 12155
rect 12759 12121 12768 12155
rect 12716 12112 12768 12121
rect 13728 12112 13780 12164
rect 11244 12044 11296 12096
rect 13360 12044 13412 12096
rect 16304 12112 16356 12164
rect 16672 12044 16724 12096
rect 2658 11942 2710 11994
rect 2722 11942 2774 11994
rect 2786 11942 2838 11994
rect 2850 11942 2902 11994
rect 2914 11942 2966 11994
rect 2978 11942 3030 11994
rect 8658 11942 8710 11994
rect 8722 11942 8774 11994
rect 8786 11942 8838 11994
rect 8850 11942 8902 11994
rect 8914 11942 8966 11994
rect 8978 11942 9030 11994
rect 14658 11942 14710 11994
rect 14722 11942 14774 11994
rect 14786 11942 14838 11994
rect 14850 11942 14902 11994
rect 14914 11942 14966 11994
rect 14978 11942 15030 11994
rect 1584 11772 1636 11824
rect 2596 11772 2648 11824
rect 2320 11636 2372 11688
rect 3056 11704 3108 11756
rect 3148 11704 3200 11756
rect 7288 11840 7340 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 8576 11840 8628 11892
rect 12440 11840 12492 11892
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 16120 11840 16172 11892
rect 12348 11772 12400 11824
rect 8300 11704 8352 11756
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 5448 11636 5500 11688
rect 8576 11636 8628 11688
rect 3700 11611 3752 11620
rect 3700 11577 3709 11611
rect 3709 11577 3743 11611
rect 3743 11577 3752 11611
rect 3700 11568 3752 11577
rect 7932 11568 7984 11620
rect 9680 11704 9732 11756
rect 10692 11704 10744 11756
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 14372 11747 14424 11756
rect 14372 11713 14381 11747
rect 14381 11713 14415 11747
rect 14415 11713 14424 11747
rect 14372 11704 14424 11713
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 14740 11636 14792 11688
rect 9588 11568 9640 11620
rect 10968 11568 11020 11620
rect 2688 11500 2740 11552
rect 8300 11500 8352 11552
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 1918 11398 1970 11450
rect 1982 11398 2034 11450
rect 2046 11398 2098 11450
rect 2110 11398 2162 11450
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 7918 11398 7970 11450
rect 7982 11398 8034 11450
rect 8046 11398 8098 11450
rect 8110 11398 8162 11450
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 13918 11398 13970 11450
rect 13982 11398 14034 11450
rect 14046 11398 14098 11450
rect 14110 11398 14162 11450
rect 14174 11398 14226 11450
rect 14238 11398 14290 11450
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 5172 11296 5224 11348
rect 10876 11296 10928 11348
rect 12072 11296 12124 11348
rect 3148 11228 3200 11280
rect 10692 11228 10744 11280
rect 12992 11296 13044 11348
rect 12900 11228 12952 11280
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 7288 11160 7340 11212
rect 8484 11160 8536 11212
rect 10416 11160 10468 11212
rect 1676 10956 1728 11008
rect 3148 10956 3200 11008
rect 3792 10956 3844 11008
rect 4068 10956 4120 11008
rect 5080 10956 5132 11008
rect 8208 11024 8260 11076
rect 9220 11092 9272 11144
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 12624 11092 12676 11144
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 17040 11228 17092 11280
rect 17224 11160 17276 11212
rect 14556 11092 14608 11144
rect 15108 11092 15160 11144
rect 16948 11092 17000 11144
rect 8484 11024 8536 11076
rect 9680 11067 9732 11076
rect 9680 11033 9689 11067
rect 9689 11033 9723 11067
rect 9723 11033 9732 11067
rect 9680 11024 9732 11033
rect 10968 11024 11020 11076
rect 12348 11024 12400 11076
rect 12716 11024 12768 11076
rect 13452 11024 13504 11076
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11244 10956 11296 10965
rect 13360 10999 13412 11008
rect 13360 10965 13369 10999
rect 13369 10965 13403 10999
rect 13403 10965 13412 10999
rect 13360 10956 13412 10965
rect 16396 10956 16448 11008
rect 2658 10854 2710 10906
rect 2722 10854 2774 10906
rect 2786 10854 2838 10906
rect 2850 10854 2902 10906
rect 2914 10854 2966 10906
rect 2978 10854 3030 10906
rect 8658 10854 8710 10906
rect 8722 10854 8774 10906
rect 8786 10854 8838 10906
rect 8850 10854 8902 10906
rect 8914 10854 8966 10906
rect 8978 10854 9030 10906
rect 14658 10854 14710 10906
rect 14722 10854 14774 10906
rect 14786 10854 14838 10906
rect 14850 10854 14902 10906
rect 14914 10854 14966 10906
rect 14978 10854 15030 10906
rect 3056 10752 3108 10804
rect 1676 10727 1728 10736
rect 1676 10693 1685 10727
rect 1685 10693 1719 10727
rect 1719 10693 1728 10727
rect 1676 10684 1728 10693
rect 4160 10752 4212 10804
rect 9680 10752 9732 10804
rect 10416 10752 10468 10804
rect 15108 10752 15160 10804
rect 3700 10684 3752 10736
rect 6460 10727 6512 10736
rect 6460 10693 6469 10727
rect 6469 10693 6503 10727
rect 6503 10693 6512 10727
rect 6460 10684 6512 10693
rect 11152 10684 11204 10736
rect 15476 10727 15528 10736
rect 10232 10659 10284 10668
rect 10232 10625 10241 10659
rect 10241 10625 10275 10659
rect 10275 10625 10284 10659
rect 10232 10616 10284 10625
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 1400 10412 1452 10464
rect 4068 10548 4120 10600
rect 15476 10693 15485 10727
rect 15485 10693 15519 10727
rect 15519 10693 15528 10727
rect 15476 10684 15528 10693
rect 15752 10727 15804 10736
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 15752 10693 15761 10727
rect 15761 10693 15795 10727
rect 15795 10693 15804 10727
rect 15752 10684 15804 10693
rect 17132 10727 17184 10736
rect 14556 10616 14608 10625
rect 14372 10548 14424 10600
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 13728 10480 13780 10532
rect 4528 10412 4580 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15108 10480 15160 10532
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 17776 10684 17828 10736
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 1918 10310 1970 10362
rect 1982 10310 2034 10362
rect 2046 10310 2098 10362
rect 2110 10310 2162 10362
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 7918 10310 7970 10362
rect 7982 10310 8034 10362
rect 8046 10310 8098 10362
rect 8110 10310 8162 10362
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 13918 10310 13970 10362
rect 13982 10310 14034 10362
rect 14046 10310 14098 10362
rect 14110 10310 14162 10362
rect 14174 10310 14226 10362
rect 14238 10310 14290 10362
rect 5540 10140 5592 10192
rect 15660 10208 15712 10260
rect 15936 10208 15988 10260
rect 4436 10004 4488 10056
rect 5356 10072 5408 10124
rect 11244 10072 11296 10124
rect 13360 10072 13412 10124
rect 14372 10115 14424 10124
rect 14372 10081 14381 10115
rect 14381 10081 14415 10115
rect 14415 10081 14424 10115
rect 14372 10072 14424 10081
rect 16396 10115 16448 10124
rect 16396 10081 16405 10115
rect 16405 10081 16439 10115
rect 16439 10081 16448 10115
rect 16396 10072 16448 10081
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 6460 10004 6512 10056
rect 10232 10004 10284 10056
rect 12624 10004 12676 10056
rect 13268 10004 13320 10056
rect 4988 9936 5040 9988
rect 5356 9936 5408 9988
rect 11428 9936 11480 9988
rect 4344 9868 4396 9920
rect 11796 9868 11848 9920
rect 13636 9868 13688 9920
rect 15384 9936 15436 9988
rect 15200 9868 15252 9920
rect 16488 9936 16540 9988
rect 16580 9868 16632 9920
rect 2658 9766 2710 9818
rect 2722 9766 2774 9818
rect 2786 9766 2838 9818
rect 2850 9766 2902 9818
rect 2914 9766 2966 9818
rect 2978 9766 3030 9818
rect 8658 9766 8710 9818
rect 8722 9766 8774 9818
rect 8786 9766 8838 9818
rect 8850 9766 8902 9818
rect 8914 9766 8966 9818
rect 8978 9766 9030 9818
rect 14658 9766 14710 9818
rect 14722 9766 14774 9818
rect 14786 9766 14838 9818
rect 14850 9766 14902 9818
rect 14914 9766 14966 9818
rect 14978 9766 15030 9818
rect 4896 9664 4948 9716
rect 5264 9664 5316 9716
rect 1768 9596 1820 9648
rect 2412 9639 2464 9648
rect 2412 9605 2421 9639
rect 2421 9605 2455 9639
rect 2455 9605 2464 9639
rect 2412 9596 2464 9605
rect 13268 9707 13320 9716
rect 13268 9673 13277 9707
rect 13277 9673 13311 9707
rect 13311 9673 13320 9707
rect 13268 9664 13320 9673
rect 10324 9596 10376 9648
rect 10876 9596 10928 9648
rect 11796 9639 11848 9648
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 12348 9596 12400 9648
rect 16764 9639 16816 9648
rect 16764 9605 16773 9639
rect 16773 9605 16807 9639
rect 16807 9605 16816 9639
rect 16764 9596 16816 9605
rect 17408 9596 17460 9648
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 3056 9528 3108 9580
rect 5080 9528 5132 9580
rect 7012 9528 7064 9580
rect 8576 9528 8628 9580
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 10692 9528 10744 9580
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 1400 9460 1452 9512
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 8484 9460 8536 9512
rect 10140 9460 10192 9512
rect 11244 9460 11296 9512
rect 12440 9460 12492 9512
rect 9220 9324 9272 9376
rect 10508 9324 10560 9376
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 1918 9222 1970 9274
rect 1982 9222 2034 9274
rect 2046 9222 2098 9274
rect 2110 9222 2162 9274
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 7918 9222 7970 9274
rect 7982 9222 8034 9274
rect 8046 9222 8098 9274
rect 8110 9222 8162 9274
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 13918 9222 13970 9274
rect 13982 9222 14034 9274
rect 14046 9222 14098 9274
rect 14110 9222 14162 9274
rect 14174 9222 14226 9274
rect 14238 9222 14290 9274
rect 6644 9120 6696 9172
rect 8576 9120 8628 9172
rect 3056 8984 3108 9036
rect 5540 8984 5592 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3700 8916 3752 8968
rect 4344 8916 4396 8968
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 7012 8916 7064 8968
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 15108 9120 15160 9172
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 5080 8848 5132 8900
rect 6000 8891 6052 8900
rect 6000 8857 6009 8891
rect 6009 8857 6043 8891
rect 6043 8857 6052 8891
rect 6000 8848 6052 8857
rect 6092 8823 6144 8832
rect 6092 8789 6101 8823
rect 6101 8789 6135 8823
rect 6135 8789 6144 8823
rect 6092 8780 6144 8789
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 7656 8916 7708 8968
rect 9220 8984 9272 9036
rect 8484 8916 8536 8968
rect 12348 9052 12400 9104
rect 10876 8984 10928 9036
rect 10692 8916 10744 8968
rect 12440 8984 12492 9036
rect 16672 8984 16724 9036
rect 17684 8984 17736 9036
rect 12348 8916 12400 8968
rect 9496 8848 9548 8900
rect 7380 8780 7432 8832
rect 10140 8780 10192 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 11428 8780 11480 8832
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 17408 8916 17460 8968
rect 13636 8891 13688 8900
rect 13636 8857 13645 8891
rect 13645 8857 13679 8891
rect 13679 8857 13688 8891
rect 13636 8848 13688 8857
rect 14372 8891 14424 8900
rect 14372 8857 14381 8891
rect 14381 8857 14415 8891
rect 14415 8857 14424 8891
rect 14372 8848 14424 8857
rect 15384 8780 15436 8832
rect 16488 8848 16540 8900
rect 16764 8848 16816 8900
rect 17132 8891 17184 8900
rect 17132 8857 17141 8891
rect 17141 8857 17175 8891
rect 17175 8857 17184 8891
rect 17132 8848 17184 8857
rect 17500 8848 17552 8900
rect 16028 8780 16080 8832
rect 16856 8780 16908 8832
rect 2658 8678 2710 8730
rect 2722 8678 2774 8730
rect 2786 8678 2838 8730
rect 2850 8678 2902 8730
rect 2914 8678 2966 8730
rect 2978 8678 3030 8730
rect 8658 8678 8710 8730
rect 8722 8678 8774 8730
rect 8786 8678 8838 8730
rect 8850 8678 8902 8730
rect 8914 8678 8966 8730
rect 8978 8678 9030 8730
rect 14658 8678 14710 8730
rect 14722 8678 14774 8730
rect 14786 8678 14838 8730
rect 14850 8678 14902 8730
rect 14914 8678 14966 8730
rect 14978 8678 15030 8730
rect 3148 8576 3200 8628
rect 3976 8576 4028 8628
rect 3056 8508 3108 8560
rect 2412 8372 2464 8424
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4528 8372 4580 8424
rect 6276 8576 6328 8628
rect 9496 8576 9548 8628
rect 10508 8619 10560 8628
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 5264 8508 5316 8560
rect 4620 8304 4672 8356
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 9956 8372 10008 8424
rect 10140 8415 10192 8424
rect 10140 8381 10149 8415
rect 10149 8381 10183 8415
rect 10183 8381 10192 8415
rect 10140 8372 10192 8381
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 7380 8304 7432 8356
rect 9772 8304 9824 8356
rect 13728 8576 13780 8628
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13452 8440 13504 8492
rect 15200 8508 15252 8560
rect 15752 8508 15804 8560
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 13728 8372 13780 8424
rect 16672 8304 16724 8356
rect 17040 8304 17092 8356
rect 2596 8236 2648 8288
rect 10416 8236 10468 8288
rect 12992 8279 13044 8288
rect 12992 8245 13001 8279
rect 13001 8245 13035 8279
rect 13035 8245 13044 8279
rect 12992 8236 13044 8245
rect 16948 8236 17000 8288
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 13918 8134 13970 8186
rect 13982 8134 14034 8186
rect 14046 8134 14098 8186
rect 14110 8134 14162 8186
rect 14174 8134 14226 8186
rect 14238 8134 14290 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 6092 8032 6144 8084
rect 7564 8032 7616 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 14372 8032 14424 8084
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 4528 7828 4580 7880
rect 5540 7760 5592 7812
rect 6828 7760 6880 7812
rect 1768 7692 1820 7744
rect 5264 7692 5316 7744
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 13820 7828 13872 7880
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 15936 7760 15988 7812
rect 16764 7760 16816 7812
rect 9220 7692 9272 7744
rect 2658 7590 2710 7642
rect 2722 7590 2774 7642
rect 2786 7590 2838 7642
rect 2850 7590 2902 7642
rect 2914 7590 2966 7642
rect 2978 7590 3030 7642
rect 8658 7590 8710 7642
rect 8722 7590 8774 7642
rect 8786 7590 8838 7642
rect 8850 7590 8902 7642
rect 8914 7590 8966 7642
rect 8978 7590 9030 7642
rect 14658 7590 14710 7642
rect 14722 7590 14774 7642
rect 14786 7590 14838 7642
rect 14850 7590 14902 7642
rect 14914 7590 14966 7642
rect 14978 7590 15030 7642
rect 1400 7284 1452 7336
rect 4804 7420 4856 7472
rect 4988 7420 5040 7472
rect 5264 7463 5316 7472
rect 5264 7429 5273 7463
rect 5273 7429 5307 7463
rect 5307 7429 5316 7463
rect 5264 7420 5316 7429
rect 6828 7488 6880 7540
rect 8576 7420 8628 7472
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 14556 7488 14608 7540
rect 9128 7420 9180 7472
rect 9404 7420 9456 7472
rect 2320 7284 2372 7336
rect 3240 7284 3292 7336
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 4804 7284 4856 7336
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10140 7352 10192 7404
rect 12440 7352 12492 7404
rect 12992 7352 13044 7404
rect 14924 7395 14976 7404
rect 14924 7361 14933 7395
rect 14933 7361 14967 7395
rect 14967 7361 14976 7395
rect 14924 7352 14976 7361
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 16580 7352 16632 7404
rect 1676 7148 1728 7200
rect 1952 7148 2004 7200
rect 3332 7148 3384 7200
rect 8668 7148 8720 7200
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 10140 7148 10192 7200
rect 12624 7148 12676 7200
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 13918 7046 13970 7098
rect 13982 7046 14034 7098
rect 14046 7046 14098 7098
rect 14110 7046 14162 7098
rect 14174 7046 14226 7098
rect 14238 7046 14290 7098
rect 9036 6944 9088 6996
rect 10140 6987 10192 6996
rect 10140 6953 10170 6987
rect 10170 6953 10192 6987
rect 10140 6944 10192 6953
rect 13820 6987 13872 6996
rect 13820 6953 13829 6987
rect 13829 6953 13863 6987
rect 13863 6953 13872 6987
rect 13820 6944 13872 6953
rect 14924 6944 14976 6996
rect 15200 6944 15252 6996
rect 16764 6944 16816 6996
rect 2320 6876 2372 6928
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 5172 6808 5224 6860
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 9404 6851 9456 6860
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 12532 6808 12584 6860
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 5540 6715 5592 6724
rect 5540 6681 5549 6715
rect 5549 6681 5583 6715
rect 5583 6681 5592 6715
rect 5540 6672 5592 6681
rect 6828 6672 6880 6724
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 8668 6740 8720 6792
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 9128 6672 9180 6724
rect 11520 6672 11572 6724
rect 11980 6715 12032 6724
rect 11980 6681 11989 6715
rect 11989 6681 12023 6715
rect 12023 6681 12032 6715
rect 11980 6672 12032 6681
rect 14096 6808 14148 6860
rect 15936 6808 15988 6860
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14372 6740 14424 6792
rect 15016 6740 15068 6792
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 12256 6604 12308 6656
rect 12348 6604 12400 6656
rect 15292 6672 15344 6724
rect 15844 6672 15896 6724
rect 14004 6604 14056 6656
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 15568 6604 15620 6613
rect 15660 6604 15712 6656
rect 16488 6672 16540 6724
rect 16856 6672 16908 6724
rect 17224 6604 17276 6656
rect 2658 6502 2710 6554
rect 2722 6502 2774 6554
rect 2786 6502 2838 6554
rect 2850 6502 2902 6554
rect 2914 6502 2966 6554
rect 2978 6502 3030 6554
rect 8658 6502 8710 6554
rect 8722 6502 8774 6554
rect 8786 6502 8838 6554
rect 8850 6502 8902 6554
rect 8914 6502 8966 6554
rect 8978 6502 9030 6554
rect 14658 6502 14710 6554
rect 14722 6502 14774 6554
rect 14786 6502 14838 6554
rect 14850 6502 14902 6554
rect 14914 6502 14966 6554
rect 14978 6502 15030 6554
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 3332 6264 3384 6316
rect 8484 6332 8536 6384
rect 12348 6400 12400 6452
rect 13820 6400 13872 6452
rect 14096 6400 14148 6452
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3792 6264 3844 6316
rect 12992 6332 13044 6384
rect 14004 6375 14056 6384
rect 14004 6341 14013 6375
rect 14013 6341 14047 6375
rect 14047 6341 14056 6375
rect 14004 6332 14056 6341
rect 15384 6400 15436 6452
rect 15292 6332 15344 6384
rect 16672 6332 16724 6384
rect 12532 6264 12584 6316
rect 15108 6264 15160 6316
rect 16856 6264 16908 6316
rect 3424 6196 3476 6205
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 3976 6128 4028 6180
rect 7564 6128 7616 6180
rect 11428 6128 11480 6180
rect 15568 6196 15620 6248
rect 2320 6060 2372 6112
rect 3884 6060 3936 6112
rect 11520 6060 11572 6112
rect 14096 6060 14148 6112
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 13918 5958 13970 6010
rect 13982 5958 14034 6010
rect 14046 5958 14098 6010
rect 14110 5958 14162 6010
rect 14174 5958 14226 6010
rect 14238 5958 14290 6010
rect 3792 5899 3844 5908
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 4620 5788 4672 5840
rect 1400 5720 1452 5772
rect 2320 5720 2372 5772
rect 3240 5720 3292 5772
rect 4068 5720 4120 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 3240 5584 3292 5636
rect 1308 5516 1360 5568
rect 1492 5516 1544 5568
rect 3332 5516 3384 5568
rect 3700 5652 3752 5704
rect 3608 5584 3660 5636
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 7012 5720 7064 5772
rect 6552 5584 6604 5636
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 8392 5720 8444 5772
rect 7656 5652 7708 5661
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 10600 5652 10652 5704
rect 11428 5788 11480 5840
rect 11152 5720 11204 5772
rect 7748 5627 7800 5636
rect 7748 5593 7757 5627
rect 7757 5593 7791 5627
rect 7791 5593 7800 5627
rect 7748 5584 7800 5593
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 12624 5720 12676 5772
rect 17224 5720 17276 5772
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 16396 5652 16448 5704
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 16764 5627 16816 5636
rect 16764 5593 16773 5627
rect 16773 5593 16807 5627
rect 16807 5593 16816 5627
rect 16764 5584 16816 5593
rect 7564 5516 7616 5568
rect 7656 5516 7708 5568
rect 11244 5516 11296 5568
rect 11428 5559 11480 5568
rect 11428 5525 11437 5559
rect 11437 5525 11471 5559
rect 11471 5525 11480 5559
rect 11428 5516 11480 5525
rect 13820 5516 13872 5568
rect 14096 5516 14148 5568
rect 15108 5516 15160 5568
rect 15292 5516 15344 5568
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 2658 5414 2710 5466
rect 2722 5414 2774 5466
rect 2786 5414 2838 5466
rect 2850 5414 2902 5466
rect 2914 5414 2966 5466
rect 2978 5414 3030 5466
rect 8658 5414 8710 5466
rect 8722 5414 8774 5466
rect 8786 5414 8838 5466
rect 8850 5414 8902 5466
rect 8914 5414 8966 5466
rect 8978 5414 9030 5466
rect 14658 5414 14710 5466
rect 14722 5414 14774 5466
rect 14786 5414 14838 5466
rect 14850 5414 14902 5466
rect 14914 5414 14966 5466
rect 14978 5414 15030 5466
rect 1400 5312 1452 5364
rect 2964 5244 3016 5296
rect 4620 5312 4672 5364
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 3700 5244 3752 5296
rect 4068 5244 4120 5296
rect 7472 5244 7524 5296
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 3608 5176 3660 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 8300 5244 8352 5296
rect 9312 5355 9364 5364
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 9312 5312 9364 5321
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 9220 5244 9272 5296
rect 14096 5312 14148 5364
rect 14372 5312 14424 5364
rect 15568 5312 15620 5364
rect 16396 5312 16448 5364
rect 13820 5287 13872 5296
rect 13820 5253 13829 5287
rect 13829 5253 13863 5287
rect 13863 5253 13872 5287
rect 13820 5244 13872 5253
rect 15108 5244 15160 5296
rect 1584 5108 1636 5160
rect 3424 5083 3476 5092
rect 3424 5049 3433 5083
rect 3433 5049 3467 5083
rect 3467 5049 3476 5083
rect 3424 5040 3476 5049
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 5172 5108 5224 5160
rect 10968 5176 11020 5228
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 5264 4972 5316 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 6828 4972 6880 5024
rect 8300 4972 8352 5024
rect 9220 4972 9272 5024
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 11336 5108 11388 5160
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16580 5244 16632 5296
rect 16764 5176 16816 5228
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 15200 5108 15252 5160
rect 17132 5151 17184 5160
rect 17132 5117 17141 5151
rect 17141 5117 17175 5151
rect 17175 5117 17184 5151
rect 17132 5108 17184 5117
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 13918 4870 13970 4922
rect 13982 4870 14034 4922
rect 14046 4870 14098 4922
rect 14110 4870 14162 4922
rect 14174 4870 14226 4922
rect 14238 4870 14290 4922
rect 7748 4768 7800 4820
rect 9680 4768 9732 4820
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 16764 4768 16816 4820
rect 17132 4768 17184 4820
rect 5172 4632 5224 4684
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 10968 4564 11020 4616
rect 15200 4632 15252 4684
rect 15936 4632 15988 4684
rect 16396 4632 16448 4684
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 16672 4564 16724 4616
rect 6828 4496 6880 4548
rect 15292 4496 15344 4548
rect 15108 4428 15160 4480
rect 2658 4326 2710 4378
rect 2722 4326 2774 4378
rect 2786 4326 2838 4378
rect 2850 4326 2902 4378
rect 2914 4326 2966 4378
rect 2978 4326 3030 4378
rect 8658 4326 8710 4378
rect 8722 4326 8774 4378
rect 8786 4326 8838 4378
rect 8850 4326 8902 4378
rect 8914 4326 8966 4378
rect 8978 4326 9030 4378
rect 14658 4326 14710 4378
rect 14722 4326 14774 4378
rect 14786 4326 14838 4378
rect 14850 4326 14902 4378
rect 14914 4326 14966 4378
rect 14978 4326 15030 4378
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 13918 3782 13970 3834
rect 13982 3782 14034 3834
rect 14046 3782 14098 3834
rect 14110 3782 14162 3834
rect 14174 3782 14226 3834
rect 14238 3782 14290 3834
rect 2658 3238 2710 3290
rect 2722 3238 2774 3290
rect 2786 3238 2838 3290
rect 2850 3238 2902 3290
rect 2914 3238 2966 3290
rect 2978 3238 3030 3290
rect 8658 3238 8710 3290
rect 8722 3238 8774 3290
rect 8786 3238 8838 3290
rect 8850 3238 8902 3290
rect 8914 3238 8966 3290
rect 8978 3238 9030 3290
rect 14658 3238 14710 3290
rect 14722 3238 14774 3290
rect 14786 3238 14838 3290
rect 14850 3238 14902 3290
rect 14914 3238 14966 3290
rect 14978 3238 15030 3290
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 13918 2694 13970 2746
rect 13982 2694 14034 2746
rect 14046 2694 14098 2746
rect 14110 2694 14162 2746
rect 14174 2694 14226 2746
rect 14238 2694 14290 2746
rect 15108 2499 15160 2508
rect 15108 2465 15117 2499
rect 15117 2465 15151 2499
rect 15151 2465 15160 2499
rect 15108 2456 15160 2465
rect 14464 2388 14516 2440
rect 2658 2150 2710 2202
rect 2722 2150 2774 2202
rect 2786 2150 2838 2202
rect 2850 2150 2902 2202
rect 2914 2150 2966 2202
rect 2978 2150 3030 2202
rect 8658 2150 8710 2202
rect 8722 2150 8774 2202
rect 8786 2150 8838 2202
rect 8850 2150 8902 2202
rect 8914 2150 8966 2202
rect 8978 2150 9030 2202
rect 14658 2150 14710 2202
rect 14722 2150 14774 2202
rect 14786 2150 14838 2202
rect 14850 2150 14902 2202
rect 14914 2150 14966 2202
rect 14978 2150 15030 2202
<< metal2 >>
rect 1122 20742 1178 21542
rect 1674 20742 1730 21542
rect 2226 20890 2282 21542
rect 2226 20862 2360 20890
rect 2226 20742 2282 20862
rect 1136 18766 1164 20742
rect 1584 18896 1636 18902
rect 1584 18838 1636 18844
rect 1124 18760 1176 18766
rect 1124 18702 1176 18708
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 16794 1440 17138
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 938 15872 994 15881
rect 938 15807 994 15816
rect 952 15502 980 15807
rect 940 15496 992 15502
rect 940 15438 992 15444
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 14822 1440 14894
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 12986 1440 14758
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 10470 1440 10542
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 9518 1440 10406
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 8974 1440 9454
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 7342 1440 8910
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 5778 1440 7278
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1308 5568 1360 5574
rect 1308 5510 1360 5516
rect 1320 5273 1348 5510
rect 1412 5370 1440 5714
rect 1504 5574 1532 18566
rect 1596 11830 1624 18838
rect 1688 18766 1716 20742
rect 1916 19068 2292 19077
rect 1972 19066 1996 19068
rect 2052 19066 2076 19068
rect 2132 19066 2156 19068
rect 2212 19066 2236 19068
rect 1972 19014 1982 19066
rect 2226 19014 2236 19066
rect 1972 19012 1996 19014
rect 2052 19012 2076 19014
rect 2132 19012 2156 19014
rect 2212 19012 2236 19014
rect 1916 19003 2292 19012
rect 2332 18766 2360 20862
rect 2778 20742 2834 21542
rect 3330 20742 3386 21542
rect 3882 20742 3938 21542
rect 4434 20890 4490 21542
rect 4434 20862 4568 20890
rect 4434 20742 4490 20862
rect 2792 18766 2820 20742
rect 3344 18766 3372 20742
rect 3896 18766 3924 20742
rect 4436 18964 4488 18970
rect 4436 18906 4488 18912
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 17882 1716 18158
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1688 14618 1716 14894
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 12918 1716 13126
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1584 11824 1636 11830
rect 1584 11766 1636 11772
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10742 1716 10950
rect 1676 10736 1728 10742
rect 1676 10678 1728 10684
rect 1780 9654 1808 18566
rect 2656 18524 3032 18533
rect 2712 18522 2736 18524
rect 2792 18522 2816 18524
rect 2872 18522 2896 18524
rect 2952 18522 2976 18524
rect 2712 18470 2722 18522
rect 2966 18470 2976 18522
rect 2712 18468 2736 18470
rect 2792 18468 2816 18470
rect 2872 18468 2896 18470
rect 2952 18468 2976 18470
rect 2656 18459 3032 18468
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2424 18222 2452 18294
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 1916 17980 2292 17989
rect 1972 17978 1996 17980
rect 2052 17978 2076 17980
rect 2132 17978 2156 17980
rect 2212 17978 2236 17980
rect 1972 17926 1982 17978
rect 2226 17926 2236 17978
rect 1972 17924 1996 17926
rect 2052 17924 2076 17926
rect 2132 17924 2156 17926
rect 2212 17924 2236 17926
rect 1916 17915 2292 17924
rect 1916 16892 2292 16901
rect 1972 16890 1996 16892
rect 2052 16890 2076 16892
rect 2132 16890 2156 16892
rect 2212 16890 2236 16892
rect 1972 16838 1982 16890
rect 2226 16838 2236 16890
rect 1972 16836 1996 16838
rect 2052 16836 2076 16838
rect 2132 16836 2156 16838
rect 2212 16836 2236 16838
rect 1916 16827 2292 16836
rect 2424 16522 2452 18158
rect 3068 17746 3096 18566
rect 3160 18426 3188 18634
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 2516 17202 2544 17682
rect 2656 17436 3032 17445
rect 2712 17434 2736 17436
rect 2792 17434 2816 17436
rect 2872 17434 2896 17436
rect 2952 17434 2976 17436
rect 2712 17382 2722 17434
rect 2966 17382 2976 17434
rect 2712 17380 2736 17382
rect 2792 17380 2816 17382
rect 2872 17380 2896 17382
rect 2952 17380 2976 17382
rect 2656 17371 3032 17380
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 3160 16658 3188 18090
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3252 17678 3280 18022
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3252 17134 3280 17478
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2656 16348 3032 16357
rect 2712 16346 2736 16348
rect 2792 16346 2816 16348
rect 2872 16346 2896 16348
rect 2952 16346 2976 16348
rect 2712 16294 2722 16346
rect 2966 16294 2976 16346
rect 2712 16292 2736 16294
rect 2792 16292 2816 16294
rect 2872 16292 2896 16294
rect 2952 16292 2976 16294
rect 2656 16283 3032 16292
rect 3160 16130 3188 16594
rect 3160 16102 3280 16130
rect 3252 16046 3280 16102
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 1916 15804 2292 15813
rect 1972 15802 1996 15804
rect 2052 15802 2076 15804
rect 2132 15802 2156 15804
rect 2212 15802 2236 15804
rect 1972 15750 1982 15802
rect 2226 15750 2236 15802
rect 1972 15748 1996 15750
rect 2052 15748 2076 15750
rect 2132 15748 2156 15750
rect 2212 15748 2236 15750
rect 1916 15739 2292 15748
rect 1916 14716 2292 14725
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 1972 14662 1982 14714
rect 2226 14662 2236 14714
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 1916 14651 2292 14660
rect 2332 14414 2360 15846
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 2656 15260 3032 15269
rect 2712 15258 2736 15260
rect 2792 15258 2816 15260
rect 2872 15258 2896 15260
rect 2952 15258 2976 15260
rect 2712 15206 2722 15258
rect 2966 15206 2976 15258
rect 2712 15204 2736 15206
rect 2792 15204 2816 15206
rect 2872 15204 2896 15206
rect 2952 15204 2976 15206
rect 2656 15195 3032 15204
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 1916 13628 2292 13637
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 1972 13574 1982 13626
rect 2226 13574 2236 13626
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 1916 13563 2292 13572
rect 2332 13326 2360 14350
rect 2424 13938 2452 14418
rect 3160 14414 3188 14758
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 14074 2544 14214
rect 2656 14172 3032 14181
rect 2712 14170 2736 14172
rect 2792 14170 2816 14172
rect 2872 14170 2896 14172
rect 2952 14170 2976 14172
rect 2712 14118 2722 14170
rect 2966 14118 2976 14170
rect 2712 14116 2736 14118
rect 2792 14116 2816 14118
rect 2872 14116 2896 14118
rect 2952 14116 2976 14118
rect 2656 14107 3032 14116
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 3160 14006 3188 14350
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 13394 2544 13670
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2656 13084 3032 13093
rect 2712 13082 2736 13084
rect 2792 13082 2816 13084
rect 2872 13082 2896 13084
rect 2952 13082 2976 13084
rect 2712 13030 2722 13082
rect 2966 13030 2976 13082
rect 2712 13028 2736 13030
rect 2792 13028 2816 13030
rect 2872 13028 2896 13030
rect 2952 13028 2976 13030
rect 2656 13019 3032 13028
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 1916 12540 2292 12549
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 1972 12486 1982 12538
rect 2226 12486 2236 12538
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 1916 12475 2292 12484
rect 2656 11996 3032 12005
rect 2712 11994 2736 11996
rect 2792 11994 2816 11996
rect 2872 11994 2896 11996
rect 2952 11994 2976 11996
rect 2712 11942 2722 11994
rect 2966 11942 2976 11994
rect 2712 11940 2736 11942
rect 2792 11940 2816 11942
rect 2872 11940 2896 11942
rect 2952 11940 2976 11942
rect 2656 11931 3032 11940
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2608 11642 2636 11766
rect 3160 11762 3188 12582
rect 3252 12170 3280 15302
rect 3436 14414 3464 18566
rect 3712 18290 3740 18566
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3804 17610 3832 18294
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 3792 17604 3844 17610
rect 3792 17546 3844 17552
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 13938 3464 14350
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 1916 11452 2292 11461
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 1972 11398 1982 11450
rect 2226 11398 2236 11450
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 1916 11387 2292 11396
rect 1916 10364 2292 10373
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 1972 10310 1982 10362
rect 2226 10310 2236 10362
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 1916 10299 2292 10308
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 2332 9586 2360 11630
rect 2608 11614 2820 11642
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2700 11150 2728 11494
rect 2792 11150 2820 11614
rect 3068 11150 3096 11698
rect 3160 11286 3188 11698
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3436 11354 3464 11630
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 2656 10908 3032 10917
rect 2712 10906 2736 10908
rect 2792 10906 2816 10908
rect 2872 10906 2896 10908
rect 2952 10906 2976 10908
rect 2712 10854 2722 10906
rect 2966 10854 2976 10906
rect 2712 10852 2736 10854
rect 2792 10852 2816 10854
rect 2872 10852 2896 10854
rect 2952 10852 2976 10854
rect 2656 10843 3032 10852
rect 3068 10810 3096 11086
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2656 9820 3032 9829
rect 2712 9818 2736 9820
rect 2792 9818 2816 9820
rect 2872 9818 2896 9820
rect 2952 9818 2976 9820
rect 2712 9766 2722 9818
rect 2966 9766 2976 9818
rect 2712 9764 2736 9766
rect 2792 9764 2816 9766
rect 2872 9764 2896 9766
rect 2952 9764 2976 9766
rect 2656 9755 3032 9764
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 1916 9276 2292 9285
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 1972 9222 1982 9274
rect 2226 9222 2236 9274
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 1916 9211 2292 9220
rect 1676 8900 1728 8906
rect 1676 8842 1728 8848
rect 1688 8090 1716 8842
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 2332 7954 2360 9318
rect 2424 8430 2452 9590
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3068 9042 3096 9522
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2656 8732 3032 8741
rect 2712 8730 2736 8732
rect 2792 8730 2816 8732
rect 2872 8730 2896 8732
rect 2952 8730 2976 8732
rect 2712 8678 2722 8730
rect 2966 8678 2976 8730
rect 2712 8676 2736 8678
rect 2792 8676 2816 8678
rect 2872 8676 2896 8678
rect 2952 8676 2976 8678
rect 2656 8667 3032 8676
rect 3068 8566 3096 8978
rect 3160 8634 3188 10950
rect 3712 10742 3740 11562
rect 3804 11014 3832 17546
rect 4356 17338 4384 18158
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4080 16250 4108 16458
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3896 15026 3924 15982
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3988 15162 4016 15302
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4080 15094 4108 16186
rect 4264 16182 4292 17002
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3896 14414 3924 14962
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 4080 13818 4108 15030
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4172 14074 4200 14894
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4080 13790 4200 13818
rect 4172 12918 4200 13790
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4172 12646 4200 12854
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 4080 10606 4108 10950
rect 4172 10810 4200 12582
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4448 10062 4476 18906
rect 4540 18766 4568 20862
rect 4986 20742 5042 21542
rect 5538 20890 5594 21542
rect 5538 20862 5672 20890
rect 5538 20742 5594 20862
rect 5000 18766 5028 20742
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5184 17678 5212 18566
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 17202 4660 17478
rect 5276 17202 5304 17750
rect 5368 17678 5396 18770
rect 5644 18766 5672 20862
rect 6090 20742 6146 21542
rect 6642 20742 6698 21542
rect 7194 20890 7250 21542
rect 7746 20890 7802 21542
rect 8298 20890 8354 21542
rect 8850 20890 8906 21542
rect 9402 20890 9458 21542
rect 9954 20890 10010 21542
rect 7194 20862 7328 20890
rect 7194 20742 7250 20862
rect 6104 18766 6132 20742
rect 6656 18766 6684 20742
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5356 17672 5408 17678
rect 5408 17620 5488 17626
rect 5356 17614 5488 17620
rect 5368 17598 5488 17614
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16590 4752 17070
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4816 16658 4844 16934
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4816 13870 4844 15438
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4816 13326 4844 13806
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12434 4844 13262
rect 4632 12406 4844 12434
rect 4632 12102 4660 12406
rect 4908 12102 4936 14214
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5000 12238 5028 13262
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3712 8974 3740 9454
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3988 8634 4016 9454
rect 4356 8974 4384 9862
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 4356 8498 4384 8910
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4540 8430 4568 10406
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2608 7886 2636 8230
rect 4540 7886 4568 8366
rect 4632 8362 4660 12038
rect 5184 11354 5212 12650
rect 5368 12646 5396 13194
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5368 12238 5396 12582
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9722 4936 9998
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5000 8498 5028 9930
rect 5092 9586 5120 10950
rect 5368 10130 5396 12038
rect 5460 11694 5488 17598
rect 5552 15570 5580 18566
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5828 17678 5856 18022
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5724 15496 5776 15502
rect 5644 15456 5724 15484
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 15162 5580 15370
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5644 14822 5672 15456
rect 5724 15438 5776 15444
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 13938 5672 14758
rect 5736 14074 5764 15302
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5920 13326 5948 18566
rect 6840 17610 6868 18838
rect 7300 18766 7328 20862
rect 7746 20862 7880 20890
rect 7746 20742 7802 20862
rect 7852 18766 7880 20862
rect 8298 20862 8432 20890
rect 8298 20742 8354 20862
rect 7916 19068 8292 19077
rect 7972 19066 7996 19068
rect 8052 19066 8076 19068
rect 8132 19066 8156 19068
rect 8212 19066 8236 19068
rect 7972 19014 7982 19066
rect 8226 19014 8236 19066
rect 7972 19012 7996 19014
rect 8052 19012 8076 19014
rect 8132 19012 8156 19014
rect 8212 19012 8236 19014
rect 7916 19003 8292 19012
rect 8404 18766 8432 20862
rect 8850 20862 8984 20890
rect 8850 20742 8906 20862
rect 8956 18766 8984 20862
rect 9402 20862 9536 20890
rect 9402 20742 9458 20862
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6932 17882 6960 18294
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6840 17270 6868 17546
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6196 15026 6224 15506
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6472 14958 6500 15302
rect 6932 15162 6960 15370
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6366 14376 6422 14385
rect 6366 14311 6368 14320
rect 6420 14311 6422 14320
rect 6368 14282 6420 14288
rect 6564 14074 6592 14962
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12986 5764 13126
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5552 12442 5580 12854
rect 5736 12850 5764 12922
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 7116 12238 7144 18566
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7208 16590 7236 17614
rect 7300 16658 7328 18362
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7300 15570 7328 16594
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7300 15026 7328 15506
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 14618 7328 14962
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7300 13394 7328 14554
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7300 12850 7328 13330
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 5448 11688 5500 11694
rect 5500 11648 5580 11676
rect 5448 11630 5500 11636
rect 5552 10198 5580 11648
rect 6472 10742 6500 12106
rect 7300 11898 7328 12786
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7300 11218 7328 11834
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5368 9994 5396 10066
rect 6472 10062 6500 10678
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 8906 5120 9522
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6798 1716 7142
rect 1780 6866 1808 7686
rect 1964 7206 1992 7822
rect 2656 7644 3032 7653
rect 2712 7642 2736 7644
rect 2792 7642 2816 7644
rect 2872 7642 2896 7644
rect 2952 7642 2976 7644
rect 2712 7590 2722 7642
rect 2966 7590 2976 7642
rect 2712 7588 2736 7590
rect 2792 7588 2816 7590
rect 2872 7588 2896 7590
rect 2952 7588 2976 7590
rect 2656 7579 3032 7588
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 2332 6934 2360 7278
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 2656 6556 3032 6565
rect 2712 6554 2736 6556
rect 2792 6554 2816 6556
rect 2872 6554 2896 6556
rect 2952 6554 2976 6556
rect 2712 6502 2722 6554
rect 2966 6502 2976 6554
rect 2712 6500 2736 6502
rect 2792 6500 2816 6502
rect 2872 6500 2896 6502
rect 2952 6500 2976 6502
rect 2656 6491 3032 6500
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 2332 5778 2360 6054
rect 3252 5778 3280 7278
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 6322 3372 7142
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1306 5264 1362 5273
rect 1306 5199 1362 5208
rect 1596 5166 1624 5646
rect 3252 5642 3280 5714
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 2656 5468 3032 5477
rect 2712 5466 2736 5468
rect 2792 5466 2816 5468
rect 2872 5466 2896 5468
rect 2952 5466 2976 5468
rect 2712 5414 2722 5466
rect 2966 5414 2976 5466
rect 2712 5412 2736 5414
rect 2792 5412 2816 5414
rect 2872 5412 2896 5414
rect 2952 5412 2976 5414
rect 2656 5403 3032 5412
rect 2964 5296 3016 5302
rect 3252 5250 3280 5578
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3016 5244 3280 5250
rect 2964 5238 3280 5244
rect 2976 5222 3280 5238
rect 3344 5234 3372 5510
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 3436 5098 3464 6190
rect 3804 5914 3832 6258
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3620 5234 3648 5578
rect 3712 5302 3740 5646
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3896 5166 3924 6054
rect 3988 5234 4016 6122
rect 4632 5846 4660 8298
rect 5092 7562 5120 8842
rect 5276 8566 5304 9658
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 9178 6684 9454
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5000 7534 5120 7562
rect 5000 7478 5028 7534
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4816 7342 4844 7414
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 5184 6866 5212 7890
rect 5552 7818 5580 8978
rect 7024 8974 7052 9522
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6012 8537 6040 8842
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5998 8528 6054 8537
rect 5998 8463 6054 8472
rect 6104 8090 6132 8774
rect 6288 8634 6316 8910
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5276 7478 5304 7686
rect 6840 7546 6868 7754
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5302 4108 5714
rect 4632 5370 4660 5782
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 5184 5166 5212 6802
rect 6840 6730 6868 7482
rect 7024 6866 7052 8910
rect 7392 8838 7420 12038
rect 7484 9058 7512 18566
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7576 17338 7604 17614
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7668 17082 7696 18566
rect 8656 18524 9032 18533
rect 8712 18522 8736 18524
rect 8792 18522 8816 18524
rect 8872 18522 8896 18524
rect 8952 18522 8976 18524
rect 8712 18470 8722 18522
rect 8966 18470 8976 18522
rect 8712 18468 8736 18470
rect 8792 18468 8816 18470
rect 8872 18468 8896 18470
rect 8952 18468 8976 18470
rect 8656 18459 9032 18468
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8220 18222 8248 18362
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 17270 7788 17682
rect 7852 17678 7880 18022
rect 7916 17980 8292 17989
rect 7972 17978 7996 17980
rect 8052 17978 8076 17980
rect 8132 17978 8156 17980
rect 8212 17978 8236 17980
rect 7972 17926 7982 17978
rect 8226 17926 8236 17978
rect 7972 17924 7996 17926
rect 8052 17924 8076 17926
rect 8132 17924 8156 17926
rect 8212 17924 8236 17926
rect 7916 17915 8292 17924
rect 8680 17882 8708 18158
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7576 17054 7696 17082
rect 7748 17128 7800 17134
rect 7852 17082 7880 17614
rect 8656 17436 9032 17445
rect 8712 17434 8736 17436
rect 8792 17434 8816 17436
rect 8872 17434 8896 17436
rect 8952 17434 8976 17436
rect 8712 17382 8722 17434
rect 8966 17382 8976 17434
rect 8712 17380 8736 17382
rect 8792 17380 8816 17382
rect 8872 17380 8896 17382
rect 8952 17380 8976 17382
rect 8656 17371 9032 17380
rect 9140 17270 9168 18294
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 7800 17076 7880 17082
rect 7748 17070 7880 17076
rect 7760 17054 7880 17070
rect 7576 12434 7604 17054
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 16658 7696 16934
rect 7916 16892 8292 16901
rect 7972 16890 7996 16892
rect 8052 16890 8076 16892
rect 8132 16890 8156 16892
rect 8212 16890 8236 16892
rect 7972 16838 7982 16890
rect 8226 16838 8236 16890
rect 7972 16836 7996 16838
rect 8052 16836 8076 16838
rect 8132 16836 8156 16838
rect 8212 16836 8236 16838
rect 7916 16827 8292 16836
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7852 15706 7880 16526
rect 8656 16348 9032 16357
rect 8712 16346 8736 16348
rect 8792 16346 8816 16348
rect 8872 16346 8896 16348
rect 8952 16346 8976 16348
rect 8712 16294 8722 16346
rect 8966 16294 8976 16346
rect 8712 16292 8736 16294
rect 8792 16292 8816 16294
rect 8872 16292 8896 16294
rect 8952 16292 8976 16294
rect 8656 16283 9032 16292
rect 7916 15804 8292 15813
rect 7972 15802 7996 15804
rect 8052 15802 8076 15804
rect 8132 15802 8156 15804
rect 8212 15802 8236 15804
rect 7972 15750 7982 15802
rect 8226 15750 8236 15802
rect 7972 15748 7996 15750
rect 8052 15748 8076 15750
rect 8132 15748 8156 15750
rect 8212 15748 8236 15750
rect 7916 15739 8292 15748
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 9140 15450 9168 17206
rect 9048 15434 9168 15450
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 9036 15428 9168 15434
rect 9088 15422 9168 15428
rect 9036 15370 9088 15376
rect 7916 14716 8292 14725
rect 7972 14714 7996 14716
rect 8052 14714 8076 14716
rect 8132 14714 8156 14716
rect 8212 14714 8236 14716
rect 7972 14662 7982 14714
rect 8226 14662 8236 14714
rect 7972 14660 7996 14662
rect 8052 14660 8076 14662
rect 8132 14660 8156 14662
rect 8212 14660 8236 14662
rect 7916 14651 8292 14660
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8128 13938 8156 14554
rect 8404 14006 8432 15370
rect 8656 15260 9032 15269
rect 8712 15258 8736 15260
rect 8792 15258 8816 15260
rect 8872 15258 8896 15260
rect 8952 15258 8976 15260
rect 8712 15206 8722 15258
rect 8966 15206 8976 15258
rect 8712 15204 8736 15206
rect 8792 15204 8816 15206
rect 8872 15204 8896 15206
rect 8952 15204 8976 15206
rect 8656 15195 9032 15204
rect 9140 15094 9168 15422
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8956 14618 8984 14894
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8758 14376 8814 14385
rect 8758 14311 8760 14320
rect 8812 14311 8814 14320
rect 8760 14282 8812 14288
rect 8656 14172 9032 14181
rect 8712 14170 8736 14172
rect 8792 14170 8816 14172
rect 8872 14170 8896 14172
rect 8952 14170 8976 14172
rect 8712 14118 8722 14170
rect 8966 14118 8976 14170
rect 8712 14116 8736 14118
rect 8792 14116 8816 14118
rect 8872 14116 8896 14118
rect 8952 14116 8976 14118
rect 8656 14107 9032 14116
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 12986 7880 13806
rect 7916 13628 8292 13637
rect 7972 13626 7996 13628
rect 8052 13626 8076 13628
rect 8132 13626 8156 13628
rect 8212 13626 8236 13628
rect 7972 13574 7982 13626
rect 8226 13574 8236 13626
rect 7972 13572 7996 13574
rect 8052 13572 8076 13574
rect 8132 13572 8156 13574
rect 8212 13572 8236 13574
rect 7916 13563 8292 13572
rect 8404 13326 8432 13942
rect 9232 13394 9260 15302
rect 9324 15162 9352 15438
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9324 14550 9352 15098
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9324 13326 9352 14350
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 8404 12986 8432 13262
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 8656 13084 9032 13093
rect 8712 13082 8736 13084
rect 8792 13082 8816 13084
rect 8872 13082 8896 13084
rect 8952 13082 8976 13084
rect 8712 13030 8722 13082
rect 8966 13030 8976 13082
rect 8712 13028 8736 13030
rect 8792 13028 8816 13030
rect 8872 13028 8896 13030
rect 8952 13028 8976 13030
rect 8656 13019 9032 13028
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 9232 12918 9260 13126
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 7916 12540 8292 12549
rect 7972 12538 7996 12540
rect 8052 12538 8076 12540
rect 8132 12538 8156 12540
rect 8212 12538 8236 12540
rect 7972 12486 7982 12538
rect 8226 12486 8236 12538
rect 7972 12484 7996 12486
rect 8052 12484 8076 12486
rect 8132 12484 8156 12486
rect 8212 12484 8236 12486
rect 7916 12475 8292 12484
rect 7576 12406 7696 12434
rect 7668 9194 7696 12406
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 7944 11626 7972 12174
rect 8128 11898 8156 12174
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8404 11762 8432 12174
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 8312 11558 8340 11698
rect 8300 11552 8352 11558
rect 8352 11512 8432 11540
rect 8300 11494 8352 11500
rect 7916 11452 8292 11461
rect 7972 11450 7996 11452
rect 8052 11450 8076 11452
rect 8132 11450 8156 11452
rect 8212 11450 8236 11452
rect 7972 11398 7982 11450
rect 8226 11398 8236 11450
rect 7972 11396 7996 11398
rect 8052 11396 8076 11398
rect 8132 11396 8156 11398
rect 8212 11396 8236 11398
rect 7916 11387 8292 11396
rect 8208 11076 8260 11082
rect 8404 11064 8432 11512
rect 8496 11218 8524 12038
rect 8588 11898 8616 12174
rect 8656 11996 9032 12005
rect 8712 11994 8736 11996
rect 8792 11994 8816 11996
rect 8872 11994 8896 11996
rect 8952 11994 8976 11996
rect 8712 11942 8722 11994
rect 8966 11942 8976 11994
rect 8712 11940 8736 11942
rect 8792 11940 8816 11942
rect 8872 11940 8896 11942
rect 8952 11940 8976 11942
rect 8656 11931 9032 11940
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8260 11036 8432 11064
rect 8484 11076 8536 11082
rect 8208 11018 8260 11024
rect 8588 11064 8616 11630
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 8536 11036 8616 11064
rect 8484 11018 8536 11024
rect 7916 10364 8292 10373
rect 7972 10362 7996 10364
rect 8052 10362 8076 10364
rect 8132 10362 8156 10364
rect 8212 10362 8236 10364
rect 7972 10310 7982 10362
rect 8226 10310 8236 10362
rect 7972 10308 7996 10310
rect 8052 10308 8076 10310
rect 8132 10308 8156 10310
rect 8212 10308 8236 10310
rect 7916 10299 8292 10308
rect 8496 9518 8524 11018
rect 8656 10908 9032 10917
rect 8712 10906 8736 10908
rect 8792 10906 8816 10908
rect 8872 10906 8896 10908
rect 8952 10906 8976 10908
rect 8712 10854 8722 10906
rect 8966 10854 8976 10906
rect 8712 10852 8736 10854
rect 8792 10852 8816 10854
rect 8872 10852 8896 10854
rect 8952 10852 8976 10854
rect 8656 10843 9032 10852
rect 8656 9820 9032 9829
rect 8712 9818 8736 9820
rect 8792 9818 8816 9820
rect 8872 9818 8896 9820
rect 8952 9818 8976 9820
rect 8712 9766 8722 9818
rect 8966 9766 8976 9818
rect 8712 9764 8736 9766
rect 8792 9764 8816 9766
rect 8872 9764 8896 9766
rect 8952 9764 8976 9766
rect 8656 9755 9032 9764
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 7916 9276 8292 9285
rect 7972 9274 7996 9276
rect 8052 9274 8076 9276
rect 8132 9274 8156 9276
rect 8212 9274 8236 9276
rect 7972 9222 7982 9274
rect 8226 9222 8236 9274
rect 7972 9220 7996 9222
rect 8052 9220 8076 9222
rect 8132 9220 8156 9222
rect 8212 9220 8236 9222
rect 7916 9211 8292 9220
rect 7668 9166 7788 9194
rect 8588 9178 8616 9522
rect 9232 9382 9260 11086
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 7484 9030 7696 9058
rect 7668 8974 7696 9030
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8362 7420 8774
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7576 8090 7604 8910
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7760 7936 7788 9166
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 7668 7908 7788 7936
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 5552 5914 5580 6666
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 5184 4690 5212 5102
rect 5276 5030 5304 5646
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6564 5166 6592 5578
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6840 5030 6868 6666
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7024 5370 7052 5714
rect 7576 5710 7604 6122
rect 7668 5710 7696 7908
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 8496 6798 8524 8910
rect 8588 7478 8616 9114
rect 9232 9042 9260 9318
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 8656 8732 9032 8741
rect 8712 8730 8736 8732
rect 8792 8730 8816 8732
rect 8872 8730 8896 8732
rect 8952 8730 8976 8732
rect 8712 8678 8722 8730
rect 8966 8678 8976 8730
rect 8712 8676 8736 8678
rect 8792 8676 8816 8678
rect 8872 8676 8896 8678
rect 8952 8676 8976 8678
rect 8656 8667 9032 8676
rect 8758 8528 8814 8537
rect 8758 8463 8814 8472
rect 8772 7886 8800 8463
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 9232 7750 9260 8978
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8656 7644 9032 7653
rect 8712 7642 8736 7644
rect 8792 7642 8816 7644
rect 8872 7642 8896 7644
rect 8952 7642 8976 7644
rect 8712 7590 8722 7642
rect 8966 7590 8976 7642
rect 8712 7588 8736 7590
rect 8792 7588 8816 7590
rect 8872 7588 8896 7590
rect 8952 7588 8976 7590
rect 8656 7579 9032 7588
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6798 8708 7142
rect 9048 7002 9076 7278
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8404 5778 8432 6598
rect 8496 6390 8524 6734
rect 9140 6730 9168 7414
rect 9232 7392 9260 7686
rect 9416 7478 9444 18838
rect 9508 18766 9536 20862
rect 9954 20862 10088 20890
rect 9954 20742 10010 20862
rect 10060 18766 10088 20862
rect 10506 20742 10562 21542
rect 11058 20742 11114 21542
rect 11610 20742 11666 21542
rect 12162 20742 12218 21542
rect 12714 20742 12770 21542
rect 13266 20890 13322 21542
rect 13266 20862 13584 20890
rect 13266 20742 13322 20862
rect 10520 18766 10548 20742
rect 11072 18766 11100 20742
rect 11624 18766 11652 20742
rect 12176 18766 12204 20742
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9784 17338 9812 17614
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9784 16590 9812 17274
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9508 14906 9536 15370
rect 9508 14878 9628 14906
rect 9600 14822 9628 14878
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9600 14482 9628 14758
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12986 9628 13126
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9600 11626 9628 12922
rect 9692 11762 9720 14826
rect 10046 14376 10102 14385
rect 10046 14311 10102 14320
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9864 11552 9916 11558
rect 10060 11540 10088 14311
rect 10152 12730 10180 18566
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 18154 10640 18226
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10244 17678 10272 18022
rect 10428 17678 10456 18022
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 16658 10272 17478
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10520 15434 10548 16390
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10612 15162 10640 18090
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10152 12702 10364 12730
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9916 11512 10088 11540
rect 9864 11494 9916 11500
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10810 9720 11018
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9508 8634 9536 8842
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9876 8537 9904 11494
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9862 8528 9918 8537
rect 9862 8463 9918 8472
rect 9968 8430 9996 9522
rect 10152 9518 10180 12174
rect 10244 10674 10272 12582
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10244 10062 10272 10610
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10336 9654 10364 12702
rect 10416 12436 10468 12442
rect 10704 12434 10732 18634
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17270 11192 17478
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16658 10916 16934
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10888 15026 10916 16594
rect 11060 16176 11112 16182
rect 10980 16124 11060 16130
rect 10980 16118 11112 16124
rect 10980 16102 11100 16118
rect 10980 15434 11008 16102
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 11060 13932 11112 13938
rect 11244 13932 11296 13938
rect 11112 13892 11192 13920
rect 11060 13874 11112 13880
rect 10416 12378 10468 12384
rect 10612 12406 10732 12434
rect 10428 11218 10456 12378
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 10810 10456 11154
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8430 10180 8774
rect 10520 8634 10548 9318
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9784 7546 9812 8298
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 10152 7410 10180 8366
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 9312 7404 9364 7410
rect 9232 7364 9312 7392
rect 9312 7346 9364 7352
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10428 7342 10456 8230
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 9416 6866 9444 7142
rect 10152 7002 10180 7142
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 8656 6556 9032 6565
rect 8712 6554 8736 6556
rect 8792 6554 8816 6556
rect 8872 6554 8896 6556
rect 8952 6554 8976 6556
rect 8712 6502 8722 6554
rect 8966 6502 8976 6554
rect 8712 6500 8736 6502
rect 8792 6500 8816 6502
rect 8872 6500 8896 6502
rect 8952 6500 8976 6502
rect 8656 6491 9032 6500
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 9324 5710 9352 6734
rect 10612 5710 10640 12406
rect 11164 12374 11192 13892
rect 11244 13874 11296 13880
rect 11256 13530 11284 13874
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11348 12306 11376 18566
rect 11612 17672 11664 17678
rect 11532 17620 11612 17626
rect 11532 17614 11664 17620
rect 11532 17598 11652 17614
rect 11532 17134 11560 17598
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11532 16046 11560 17070
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11716 15094 11744 18566
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 17746 12112 18022
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11808 15570 11836 15846
rect 11900 15706 11928 15982
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11808 15026 11836 15506
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 14346 11836 14962
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10704 11286 10732 11698
rect 10888 11354 10916 12174
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10980 11082 11008 11562
rect 11256 11150 11284 12038
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11244 11144 11296 11150
rect 11164 11104 11244 11132
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 11164 10742 11192 11104
rect 11348 11121 11376 11698
rect 11244 11086 11296 11092
rect 11334 11112 11390 11121
rect 11334 11047 11390 11056
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11256 10130 11284 10950
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11440 9994 11468 13942
rect 11808 13308 11836 14282
rect 12176 14006 12204 18566
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12268 17542 12296 18158
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12452 16574 12480 18906
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12452 16546 12572 16574
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 11888 13320 11940 13326
rect 11808 13280 11888 13308
rect 11808 11762 11836 13280
rect 11888 13262 11940 13268
rect 11992 13138 12020 13670
rect 12176 13394 12204 13670
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12072 13184 12124 13190
rect 11992 13132 12072 13138
rect 11992 13126 12124 13132
rect 11992 13110 12112 13126
rect 11992 12850 12020 13110
rect 12176 12850 12204 13330
rect 12360 12986 12388 13330
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12452 11898 12480 12854
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12084 11354 12112 11630
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12360 11082 12388 11766
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10704 9178 10732 9522
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10704 8974 10732 9114
rect 10888 9042 10916 9590
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8498 10824 8774
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 7576 5574 7604 5646
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 5386 7696 5510
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7484 5358 7696 5386
rect 7484 5302 7512 5358
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6380 4690 6408 4966
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6840 4554 6868 4966
rect 7760 4826 7788 5578
rect 8656 5468 9032 5477
rect 8712 5466 8736 5468
rect 8792 5466 8816 5468
rect 8872 5466 8896 5468
rect 8952 5466 8976 5468
rect 8712 5414 8722 5466
rect 8966 5414 8976 5466
rect 8712 5412 8736 5414
rect 8792 5412 8816 5414
rect 8872 5412 8896 5414
rect 8952 5412 8976 5414
rect 8656 5403 9032 5412
rect 9324 5370 9352 5646
rect 11164 5370 11192 5714
rect 11256 5710 11284 9454
rect 11440 8838 11468 9930
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11808 9654 11836 9862
rect 12360 9654 12388 11018
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12360 9110 12388 9590
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12360 8974 12388 9046
rect 12452 9042 12480 9454
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11440 6186 11468 8774
rect 12452 8090 12480 8978
rect 12544 8498 12572 16546
rect 12636 12238 12664 18838
rect 12728 18766 12756 20742
rect 13556 18766 13584 20862
rect 13818 20742 13874 21542
rect 14370 20890 14426 21542
rect 14922 20890 14978 21542
rect 15474 20890 15530 21542
rect 16026 20890 16082 21542
rect 16578 20890 16634 21542
rect 17130 20890 17186 21542
rect 14370 20862 14504 20890
rect 14370 20742 14426 20862
rect 13832 18766 13860 20742
rect 13916 19068 14292 19077
rect 13972 19066 13996 19068
rect 14052 19066 14076 19068
rect 14132 19066 14156 19068
rect 14212 19066 14236 19068
rect 13972 19014 13982 19066
rect 14226 19014 14236 19066
rect 13972 19012 13996 19014
rect 14052 19012 14076 19014
rect 14132 19012 14156 19014
rect 14212 19012 14236 19014
rect 13916 19003 14292 19012
rect 14476 18766 14504 20862
rect 14922 20862 15056 20890
rect 14922 20742 14978 20862
rect 15028 18766 15056 20862
rect 15474 20862 15608 20890
rect 15474 20742 15530 20862
rect 15580 18766 15608 20862
rect 16026 20862 16344 20890
rect 16026 20742 16082 20862
rect 16316 18766 16344 20862
rect 16578 20862 16896 20890
rect 16578 20742 16634 20862
rect 16868 18766 16896 20862
rect 17130 20862 17264 20890
rect 17130 20742 17186 20862
rect 17236 18766 17264 20862
rect 17682 20742 17738 21542
rect 18234 20742 18290 21542
rect 17696 18766 17724 20742
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17882 12848 18022
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 13004 16574 13032 18566
rect 13372 18426 13400 18566
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13464 18306 13492 18362
rect 13740 18358 13768 18566
rect 13372 18290 13492 18306
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 14568 18290 14596 18566
rect 14656 18524 15032 18533
rect 14712 18522 14736 18524
rect 14792 18522 14816 18524
rect 14872 18522 14896 18524
rect 14952 18522 14976 18524
rect 14712 18470 14722 18522
rect 14966 18470 14976 18522
rect 14712 18468 14736 18470
rect 14792 18468 14816 18470
rect 14872 18468 14896 18470
rect 14952 18468 14976 18470
rect 14656 18459 15032 18468
rect 13360 18284 13492 18290
rect 13412 18278 13492 18284
rect 13544 18284 13596 18290
rect 13360 18226 13412 18232
rect 13544 18226 13596 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 13084 16584 13136 16590
rect 13004 16546 13084 16574
rect 13372 16574 13400 18226
rect 13556 17882 13584 18226
rect 13916 17980 14292 17989
rect 13972 17978 13996 17980
rect 14052 17978 14076 17980
rect 14132 17978 14156 17980
rect 14212 17978 14236 17980
rect 13972 17926 13982 17978
rect 14226 17926 14236 17978
rect 13972 17924 13996 17926
rect 14052 17924 14076 17926
rect 14132 17924 14156 17926
rect 14212 17924 14236 17926
rect 13916 17915 14292 17924
rect 15212 17882 15240 18226
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13372 16546 13492 16574
rect 13084 16526 13136 16532
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12728 15638 12756 16390
rect 13096 16114 13124 16526
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13280 16182 13308 16458
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 13280 16046 13308 16118
rect 13464 16114 13492 16546
rect 13832 16454 13860 17546
rect 13916 16892 14292 16901
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14156 16892
rect 14212 16890 14236 16892
rect 13972 16838 13982 16890
rect 14226 16838 14236 16890
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14156 16838
rect 14212 16836 14236 16838
rect 13916 16827 14292 16836
rect 14568 16658 14596 17682
rect 14656 17436 15032 17445
rect 14712 17434 14736 17436
rect 14792 17434 14816 17436
rect 14872 17434 14896 17436
rect 14952 17434 14976 17436
rect 14712 17382 14722 17434
rect 14966 17382 14976 17434
rect 14712 17380 14736 17382
rect 14792 17380 14816 17382
rect 14872 17380 14896 17382
rect 14952 17380 14976 17382
rect 14656 17371 15032 17380
rect 15304 17202 15332 18022
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16250 13860 16390
rect 14200 16250 14228 16458
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 12728 15502 12756 15574
rect 13464 15502 13492 15574
rect 13648 15502 13676 15846
rect 13916 15804 14292 15813
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14156 15804
rect 14212 15802 14236 15804
rect 13972 15750 13982 15802
rect 14226 15750 14236 15802
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14156 15750
rect 14212 15748 14236 15750
rect 13916 15739 14292 15748
rect 14568 15586 14596 16594
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 14656 16348 15032 16357
rect 14712 16346 14736 16348
rect 14792 16346 14816 16348
rect 14872 16346 14896 16348
rect 14952 16346 14976 16348
rect 14712 16294 14722 16346
rect 14966 16294 14976 16346
rect 14712 16292 14736 16294
rect 14792 16292 14816 16294
rect 14872 16292 14896 16294
rect 14952 16292 14976 16294
rect 14656 16283 15032 16292
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14752 15706 14780 15982
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14476 15558 14596 15586
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12636 11234 12664 12174
rect 12728 12170 12756 15098
rect 13542 14376 13598 14385
rect 13542 14311 13544 14320
rect 13596 14311 13598 14320
rect 13544 14282 13596 14288
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12986 12848 13262
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 13832 12782 13860 15302
rect 14384 15162 14412 15370
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 13916 14716 14292 14725
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14156 14716
rect 14212 14714 14236 14716
rect 13972 14662 13982 14714
rect 14226 14662 14236 14714
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14156 14662
rect 14212 14660 14236 14662
rect 13916 14651 14292 14660
rect 14384 14346 14412 14758
rect 14476 14482 14504 15558
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 14958 14596 15438
rect 14656 15260 15032 15269
rect 14712 15258 14736 15260
rect 14792 15258 14816 15260
rect 14872 15258 14896 15260
rect 14952 15258 14976 15260
rect 14712 15206 14722 15258
rect 14966 15206 14976 15258
rect 14712 15204 14736 15206
rect 14792 15204 14816 15206
rect 14872 15204 14896 15206
rect 14952 15204 14976 15206
rect 14656 15195 15032 15204
rect 15120 15026 15148 16050
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14476 14006 14504 14418
rect 14656 14172 15032 14181
rect 14712 14170 14736 14172
rect 14792 14170 14816 14172
rect 14872 14170 14896 14172
rect 14952 14170 14976 14172
rect 14712 14118 14722 14170
rect 14966 14118 14976 14170
rect 14712 14116 14736 14118
rect 14792 14116 14816 14118
rect 14872 14116 14896 14118
rect 14952 14116 14976 14118
rect 14656 14107 15032 14116
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 13916 13628 14292 13637
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14156 13628
rect 14212 13626 14236 13628
rect 13972 13574 13982 13626
rect 14226 13574 14236 13626
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14156 13574
rect 14212 13572 14236 13574
rect 13916 13563 14292 13572
rect 14476 12832 14504 13942
rect 14656 13084 15032 13093
rect 14712 13082 14736 13084
rect 14792 13082 14816 13084
rect 14872 13082 14896 13084
rect 14952 13082 14976 13084
rect 14712 13030 14722 13082
rect 14966 13030 14976 13082
rect 14712 13028 14736 13030
rect 14792 13028 14816 13030
rect 14872 13028 14896 13030
rect 14952 13028 14976 13030
rect 14656 13019 15032 13028
rect 14556 12844 14608 12850
rect 14476 12804 14556 12832
rect 14556 12786 14608 12792
rect 15120 12782 15148 14962
rect 15304 14498 15332 16390
rect 15396 14890 15424 18158
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15488 17338 15516 17546
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15488 15026 15516 15914
rect 15580 15026 15608 18566
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15672 17270 15700 18022
rect 15660 17264 15712 17270
rect 15660 17206 15712 17212
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15304 14470 15424 14498
rect 15396 14346 15424 14470
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15396 13258 15424 14282
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15396 12918 15424 13194
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 13916 12540 14292 12549
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14156 12540
rect 14212 12538 14236 12540
rect 13972 12486 13982 12538
rect 14226 12486 14236 12538
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14156 12486
rect 14212 12484 14236 12486
rect 13916 12475 14292 12484
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12900 11280 12952 11286
rect 12636 11206 12756 11234
rect 12900 11222 12952 11228
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12636 10062 12664 11086
rect 12728 11082 12756 11206
rect 12912 11150 12940 11222
rect 13004 11150 13032 11290
rect 13372 11150 13400 12038
rect 13556 11898 13584 12174
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13360 11144 13412 11150
rect 13556 11098 13584 11834
rect 13360 11086 13412 11092
rect 13464 11082 13584 11098
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 13452 11076 13584 11082
rect 13504 11070 13584 11076
rect 13452 11018 13504 11024
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10130 13400 10950
rect 13740 10538 13768 12106
rect 14656 11996 15032 12005
rect 14712 11994 14736 11996
rect 14792 11994 14816 11996
rect 14872 11994 14896 11996
rect 14952 11994 14976 11996
rect 14712 11942 14722 11994
rect 14966 11942 14976 11994
rect 14712 11940 14736 11942
rect 14792 11940 14816 11942
rect 14872 11940 14896 11942
rect 14952 11940 14976 11942
rect 14656 11931 15032 11940
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 13916 11452 14292 11461
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14156 11452
rect 14212 11450 14236 11452
rect 13972 11398 13982 11450
rect 14226 11398 14236 11450
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14156 11398
rect 14212 11396 14236 11398
rect 13916 11387 14292 11396
rect 14384 10606 14412 11698
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14752 11354 14780 11630
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 14568 10674 14596 11086
rect 14656 10908 15032 10917
rect 14712 10906 14736 10908
rect 14792 10906 14816 10908
rect 14872 10906 14896 10908
rect 14952 10906 14976 10908
rect 14712 10854 14722 10906
rect 14966 10854 14976 10906
rect 14712 10852 14736 10854
rect 14792 10852 14816 10854
rect 14872 10852 14896 10854
rect 14952 10852 14976 10854
rect 14656 10843 15032 10852
rect 15120 10810 15148 11086
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15488 10742 15516 14962
rect 15672 14890 15700 14962
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15672 10674 15700 14826
rect 15764 10742 15792 18566
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13280 9722 13308 9998
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13648 8906 13676 9862
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13740 8634 13768 10474
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 13916 10364 14292 10373
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14156 10364
rect 14212 10362 14236 10364
rect 13972 10310 13982 10362
rect 14226 10310 14236 10362
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14156 10310
rect 14212 10308 14236 10310
rect 13916 10299 14292 10308
rect 14384 10130 14412 10406
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14656 9820 15032 9829
rect 14712 9818 14736 9820
rect 14792 9818 14816 9820
rect 14872 9818 14896 9820
rect 14952 9818 14976 9820
rect 14712 9766 14722 9818
rect 14966 9766 14976 9818
rect 14712 9764 14736 9766
rect 14792 9764 14816 9766
rect 14872 9764 14896 9766
rect 14952 9764 14976 9766
rect 14656 9755 15032 9764
rect 13916 9276 14292 9285
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14156 9276
rect 14212 9274 14236 9276
rect 13972 9222 13982 9274
rect 14226 9222 14236 9274
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14156 9222
rect 14212 9220 14236 9222
rect 13916 9211 14292 9220
rect 15120 9178 15148 10474
rect 15672 10266 15700 10610
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13818 8528 13874 8537
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 13452 8492 13504 8498
rect 13818 8463 13874 8472
rect 13452 8434 13504 8440
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12452 7410 12480 8026
rect 13004 7410 13032 8230
rect 12440 7404 12492 7410
rect 12992 7404 13044 7410
rect 12492 7364 12572 7392
rect 12440 7346 12492 7352
rect 12544 6866 12572 7364
rect 12992 7346 13044 7352
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11440 5846 11468 6122
rect 11532 6118 11560 6666
rect 11992 6458 12020 6666
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 12268 6254 12296 6598
rect 12360 6458 12388 6598
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12544 6322 12572 6802
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 12268 5710 12296 6190
rect 12636 5778 12664 7142
rect 13004 6390 13032 7346
rect 13464 6866 13492 8434
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13740 6798 13768 8366
rect 13832 7886 13860 8463
rect 13916 8188 14292 8197
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14156 8188
rect 14212 8186 14236 8188
rect 13972 8134 13982 8186
rect 14226 8134 14236 8186
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14156 8134
rect 14212 8132 14236 8134
rect 13916 8123 14292 8132
rect 14384 8090 14412 8842
rect 14656 8732 15032 8741
rect 14712 8730 14736 8732
rect 14792 8730 14816 8732
rect 14872 8730 14896 8732
rect 14952 8730 14976 8732
rect 14712 8678 14722 8730
rect 14966 8678 14976 8730
rect 14712 8676 14736 8678
rect 14792 8676 14816 8678
rect 14872 8676 14896 8678
rect 14952 8676 14976 8678
rect 14656 8667 15032 8676
rect 15212 8566 15240 9862
rect 15396 8838 15424 9930
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15200 8560 15252 8566
rect 14646 8528 14702 8537
rect 15200 8502 15252 8508
rect 14646 8463 14648 8472
rect 14700 8463 14702 8472
rect 14648 8434 14700 8440
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 13916 7100 14292 7109
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14156 7100
rect 14212 7098 14236 7100
rect 13972 7046 13982 7098
rect 14226 7046 14236 7098
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14156 7046
rect 14212 7044 14236 7046
rect 13916 7035 14292 7044
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13832 6458 13860 6938
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14016 6390 14044 6598
rect 14108 6458 14136 6802
rect 14372 6792 14424 6798
rect 14476 6746 14504 7822
rect 14568 7546 14596 7890
rect 14656 7644 15032 7653
rect 14712 7642 14736 7644
rect 14792 7642 14816 7644
rect 14872 7642 14896 7644
rect 14952 7642 14976 7644
rect 14712 7590 14722 7642
rect 14966 7590 14976 7642
rect 14712 7588 14736 7590
rect 14792 7588 14816 7590
rect 14872 7588 14896 7590
rect 14952 7588 14976 7590
rect 14656 7579 15032 7588
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 14936 7002 14964 7346
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 15028 6798 15056 7346
rect 15212 7002 15240 7346
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 14424 6740 14504 6746
rect 14372 6734 14504 6740
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 14384 6718 14504 6734
rect 15292 6724 15344 6730
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14108 6118 14136 6394
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13916 6012 14292 6021
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14156 6012
rect 14212 6010 14236 6012
rect 13972 5958 13982 6010
rect 14226 5958 14236 6010
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14156 5958
rect 14212 5956 14236 5958
rect 13916 5947 14292 5956
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 8312 5030 8340 5238
rect 9232 5030 9260 5238
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 9692 4826 9720 5102
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 10980 4622 11008 5170
rect 11256 4622 11284 5510
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11348 4826 11376 5102
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11440 4622 11468 5510
rect 13832 5302 13860 5510
rect 14108 5370 14136 5510
rect 14384 5370 14412 6718
rect 15292 6666 15344 6672
rect 14656 6556 15032 6565
rect 14712 6554 14736 6556
rect 14792 6554 14816 6556
rect 14872 6554 14896 6556
rect 14952 6554 14976 6556
rect 14712 6502 14722 6554
rect 14966 6502 14976 6554
rect 14712 6500 14736 6502
rect 14792 6500 14816 6502
rect 14872 6500 14896 6502
rect 14952 6500 14976 6502
rect 14656 6491 15032 6500
rect 15304 6390 15332 6666
rect 15396 6458 15424 6734
rect 15672 6662 15700 10202
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15764 7954 15792 8502
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15856 6730 15884 18566
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 15948 18086 15976 18226
rect 16132 18154 16160 18226
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 16224 17134 16252 18226
rect 16684 18057 16712 18566
rect 16670 18048 16726 18057
rect 16670 17983 16726 17992
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16224 16794 16252 17070
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16316 16522 16344 17546
rect 17328 16574 17356 18566
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17604 17610 17632 18090
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17328 16546 17448 16574
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 16250 16160 16390
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16132 15502 16160 16186
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15948 14618 15976 14962
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 11898 16160 12718
rect 16316 12170 16344 13194
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16592 12306 16620 12786
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16684 12102 16712 12582
rect 16776 12442 16804 16118
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17052 15502 17080 15846
rect 17328 15502 17356 15846
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 17052 13870 17080 15302
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 12782 16988 13126
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10266 15976 10610
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16408 10130 16436 10950
rect 16776 10674 16804 12378
rect 16960 11150 16988 12718
rect 17052 11286 17080 13806
rect 17144 13734 17172 13874
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 12782 17172 13670
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16500 8906 16528 9930
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 8974 16620 9862
rect 16776 9654 16804 10610
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 17052 9382 17080 11222
rect 17236 11218 17264 13806
rect 17328 12986 17356 13874
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16040 7954 16068 8774
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15948 6866 15976 7754
rect 16592 7410 16620 8910
rect 16684 8498 16712 8978
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5574 15148 6258
rect 15580 6254 15608 6598
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 14656 5468 15032 5477
rect 14712 5466 14736 5468
rect 14792 5466 14816 5468
rect 14872 5466 14896 5468
rect 14952 5466 14976 5468
rect 14712 5414 14722 5466
rect 14966 5414 14976 5466
rect 14712 5412 14736 5414
rect 14792 5412 14816 5414
rect 14872 5412 14896 5414
rect 14952 5412 14976 5414
rect 14656 5403 15032 5412
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 15120 5302 15148 5510
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 13916 4924 14292 4933
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14156 4924
rect 14212 4922 14236 4924
rect 13972 4870 13982 4922
rect 14226 4870 14236 4922
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14156 4870
rect 14212 4868 14236 4870
rect 13916 4859 14292 4868
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 15120 4486 15148 5238
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15212 4690 15240 5102
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15304 4554 15332 5510
rect 15580 5370 15608 6190
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15948 5234 15976 6802
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16500 5710 16528 6666
rect 16684 6390 16712 8298
rect 16776 7818 16804 8842
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 8498 16896 8774
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 17052 8362 17080 9318
rect 17144 8906 17172 10678
rect 17420 9654 17448 16546
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17604 15910 17632 16458
rect 17696 16182 17724 18022
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17512 12850 17540 13942
rect 17604 13394 17632 15302
rect 17788 14074 17816 18566
rect 18248 18290 18276 20742
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 16658 17908 17682
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 14482 17908 16594
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17788 13274 17816 14010
rect 17880 13394 17908 14418
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17788 13246 17908 13274
rect 17880 12850 17908 13246
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17512 12442 17540 12786
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17788 10742 17816 12786
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17420 8974 17448 9590
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17512 8906 17540 9522
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 9042 17724 9318
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16776 7698 16804 7754
rect 16776 7670 16896 7698
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 7002 16804 7142
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16868 6730 16896 7670
rect 16960 7342 16988 8230
rect 17512 8090 17540 8842
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16868 6322 16896 6666
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16578 5808 16634 5817
rect 17236 5778 17264 6598
rect 16578 5743 16634 5752
rect 17224 5772 17276 5778
rect 16592 5710 16620 5743
rect 17224 5714 17276 5720
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16408 5370 16436 5646
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15948 4690 15976 5170
rect 16408 4690 16436 5306
rect 16592 5302 16620 5646
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16684 4622 16712 5510
rect 16776 5234 16804 5578
rect 17236 5234 17264 5714
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 16776 4826 16804 5170
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17144 4826 17172 5102
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 2656 4380 3032 4389
rect 2712 4378 2736 4380
rect 2792 4378 2816 4380
rect 2872 4378 2896 4380
rect 2952 4378 2976 4380
rect 2712 4326 2722 4378
rect 2966 4326 2976 4378
rect 2712 4324 2736 4326
rect 2792 4324 2816 4326
rect 2872 4324 2896 4326
rect 2952 4324 2976 4326
rect 2656 4315 3032 4324
rect 8656 4380 9032 4389
rect 8712 4378 8736 4380
rect 8792 4378 8816 4380
rect 8872 4378 8896 4380
rect 8952 4378 8976 4380
rect 8712 4326 8722 4378
rect 8966 4326 8976 4378
rect 8712 4324 8736 4326
rect 8792 4324 8816 4326
rect 8872 4324 8896 4326
rect 8952 4324 8976 4326
rect 8656 4315 9032 4324
rect 14656 4380 15032 4389
rect 14712 4378 14736 4380
rect 14792 4378 14816 4380
rect 14872 4378 14896 4380
rect 14952 4378 14976 4380
rect 14712 4326 14722 4378
rect 14966 4326 14976 4378
rect 14712 4324 14736 4326
rect 14792 4324 14816 4326
rect 14872 4324 14896 4326
rect 14952 4324 14976 4326
rect 14656 4315 15032 4324
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 13916 3836 14292 3845
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14156 3836
rect 14212 3834 14236 3836
rect 13972 3782 13982 3834
rect 14226 3782 14236 3834
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14156 3782
rect 14212 3780 14236 3782
rect 13916 3771 14292 3780
rect 2656 3292 3032 3301
rect 2712 3290 2736 3292
rect 2792 3290 2816 3292
rect 2872 3290 2896 3292
rect 2952 3290 2976 3292
rect 2712 3238 2722 3290
rect 2966 3238 2976 3290
rect 2712 3236 2736 3238
rect 2792 3236 2816 3238
rect 2872 3236 2896 3238
rect 2952 3236 2976 3238
rect 2656 3227 3032 3236
rect 8656 3292 9032 3301
rect 8712 3290 8736 3292
rect 8792 3290 8816 3292
rect 8872 3290 8896 3292
rect 8952 3290 8976 3292
rect 8712 3238 8722 3290
rect 8966 3238 8976 3290
rect 8712 3236 8736 3238
rect 8792 3236 8816 3238
rect 8872 3236 8896 3238
rect 8952 3236 8976 3238
rect 8656 3227 9032 3236
rect 14656 3292 15032 3301
rect 14712 3290 14736 3292
rect 14792 3290 14816 3292
rect 14872 3290 14896 3292
rect 14952 3290 14976 3292
rect 14712 3238 14722 3290
rect 14966 3238 14976 3290
rect 14712 3236 14736 3238
rect 14792 3236 14816 3238
rect 14872 3236 14896 3238
rect 14952 3236 14976 3238
rect 14656 3227 15032 3236
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 13916 2748 14292 2757
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14156 2748
rect 14212 2746 14236 2748
rect 13972 2694 13982 2746
rect 14226 2694 14236 2746
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14156 2694
rect 14212 2692 14236 2694
rect 13916 2683 14292 2692
rect 15120 2514 15148 4422
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 2656 2204 3032 2213
rect 2712 2202 2736 2204
rect 2792 2202 2816 2204
rect 2872 2202 2896 2204
rect 2952 2202 2976 2204
rect 2712 2150 2722 2202
rect 2966 2150 2976 2202
rect 2712 2148 2736 2150
rect 2792 2148 2816 2150
rect 2872 2148 2896 2150
rect 2952 2148 2976 2150
rect 2656 2139 3032 2148
rect 8656 2204 9032 2213
rect 8712 2202 8736 2204
rect 8792 2202 8816 2204
rect 8872 2202 8896 2204
rect 8952 2202 8976 2204
rect 8712 2150 8722 2202
rect 8966 2150 8976 2202
rect 8712 2148 8736 2150
rect 8792 2148 8816 2150
rect 8872 2148 8896 2150
rect 8952 2148 8976 2150
rect 8656 2139 9032 2148
rect 14476 800 14504 2382
rect 14656 2204 15032 2213
rect 14712 2202 14736 2204
rect 14792 2202 14816 2204
rect 14872 2202 14896 2204
rect 14952 2202 14976 2204
rect 14712 2150 14722 2202
rect 14966 2150 14976 2202
rect 14712 2148 14736 2150
rect 14792 2148 14816 2150
rect 14872 2148 14896 2150
rect 14952 2148 14976 2150
rect 14656 2139 15032 2148
rect 14462 0 14518 800
<< via2 >>
rect 938 15816 994 15872
rect 1916 19066 1972 19068
rect 1996 19066 2052 19068
rect 2076 19066 2132 19068
rect 2156 19066 2212 19068
rect 2236 19066 2292 19068
rect 1916 19014 1918 19066
rect 1918 19014 1970 19066
rect 1970 19014 1972 19066
rect 1996 19014 2034 19066
rect 2034 19014 2046 19066
rect 2046 19014 2052 19066
rect 2076 19014 2098 19066
rect 2098 19014 2110 19066
rect 2110 19014 2132 19066
rect 2156 19014 2162 19066
rect 2162 19014 2174 19066
rect 2174 19014 2212 19066
rect 2236 19014 2238 19066
rect 2238 19014 2290 19066
rect 2290 19014 2292 19066
rect 1916 19012 1972 19014
rect 1996 19012 2052 19014
rect 2076 19012 2132 19014
rect 2156 19012 2212 19014
rect 2236 19012 2292 19014
rect 2656 18522 2712 18524
rect 2736 18522 2792 18524
rect 2816 18522 2872 18524
rect 2896 18522 2952 18524
rect 2976 18522 3032 18524
rect 2656 18470 2658 18522
rect 2658 18470 2710 18522
rect 2710 18470 2712 18522
rect 2736 18470 2774 18522
rect 2774 18470 2786 18522
rect 2786 18470 2792 18522
rect 2816 18470 2838 18522
rect 2838 18470 2850 18522
rect 2850 18470 2872 18522
rect 2896 18470 2902 18522
rect 2902 18470 2914 18522
rect 2914 18470 2952 18522
rect 2976 18470 2978 18522
rect 2978 18470 3030 18522
rect 3030 18470 3032 18522
rect 2656 18468 2712 18470
rect 2736 18468 2792 18470
rect 2816 18468 2872 18470
rect 2896 18468 2952 18470
rect 2976 18468 3032 18470
rect 1916 17978 1972 17980
rect 1996 17978 2052 17980
rect 2076 17978 2132 17980
rect 2156 17978 2212 17980
rect 2236 17978 2292 17980
rect 1916 17926 1918 17978
rect 1918 17926 1970 17978
rect 1970 17926 1972 17978
rect 1996 17926 2034 17978
rect 2034 17926 2046 17978
rect 2046 17926 2052 17978
rect 2076 17926 2098 17978
rect 2098 17926 2110 17978
rect 2110 17926 2132 17978
rect 2156 17926 2162 17978
rect 2162 17926 2174 17978
rect 2174 17926 2212 17978
rect 2236 17926 2238 17978
rect 2238 17926 2290 17978
rect 2290 17926 2292 17978
rect 1916 17924 1972 17926
rect 1996 17924 2052 17926
rect 2076 17924 2132 17926
rect 2156 17924 2212 17926
rect 2236 17924 2292 17926
rect 1916 16890 1972 16892
rect 1996 16890 2052 16892
rect 2076 16890 2132 16892
rect 2156 16890 2212 16892
rect 2236 16890 2292 16892
rect 1916 16838 1918 16890
rect 1918 16838 1970 16890
rect 1970 16838 1972 16890
rect 1996 16838 2034 16890
rect 2034 16838 2046 16890
rect 2046 16838 2052 16890
rect 2076 16838 2098 16890
rect 2098 16838 2110 16890
rect 2110 16838 2132 16890
rect 2156 16838 2162 16890
rect 2162 16838 2174 16890
rect 2174 16838 2212 16890
rect 2236 16838 2238 16890
rect 2238 16838 2290 16890
rect 2290 16838 2292 16890
rect 1916 16836 1972 16838
rect 1996 16836 2052 16838
rect 2076 16836 2132 16838
rect 2156 16836 2212 16838
rect 2236 16836 2292 16838
rect 2656 17434 2712 17436
rect 2736 17434 2792 17436
rect 2816 17434 2872 17436
rect 2896 17434 2952 17436
rect 2976 17434 3032 17436
rect 2656 17382 2658 17434
rect 2658 17382 2710 17434
rect 2710 17382 2712 17434
rect 2736 17382 2774 17434
rect 2774 17382 2786 17434
rect 2786 17382 2792 17434
rect 2816 17382 2838 17434
rect 2838 17382 2850 17434
rect 2850 17382 2872 17434
rect 2896 17382 2902 17434
rect 2902 17382 2914 17434
rect 2914 17382 2952 17434
rect 2976 17382 2978 17434
rect 2978 17382 3030 17434
rect 3030 17382 3032 17434
rect 2656 17380 2712 17382
rect 2736 17380 2792 17382
rect 2816 17380 2872 17382
rect 2896 17380 2952 17382
rect 2976 17380 3032 17382
rect 2656 16346 2712 16348
rect 2736 16346 2792 16348
rect 2816 16346 2872 16348
rect 2896 16346 2952 16348
rect 2976 16346 3032 16348
rect 2656 16294 2658 16346
rect 2658 16294 2710 16346
rect 2710 16294 2712 16346
rect 2736 16294 2774 16346
rect 2774 16294 2786 16346
rect 2786 16294 2792 16346
rect 2816 16294 2838 16346
rect 2838 16294 2850 16346
rect 2850 16294 2872 16346
rect 2896 16294 2902 16346
rect 2902 16294 2914 16346
rect 2914 16294 2952 16346
rect 2976 16294 2978 16346
rect 2978 16294 3030 16346
rect 3030 16294 3032 16346
rect 2656 16292 2712 16294
rect 2736 16292 2792 16294
rect 2816 16292 2872 16294
rect 2896 16292 2952 16294
rect 2976 16292 3032 16294
rect 1916 15802 1972 15804
rect 1996 15802 2052 15804
rect 2076 15802 2132 15804
rect 2156 15802 2212 15804
rect 2236 15802 2292 15804
rect 1916 15750 1918 15802
rect 1918 15750 1970 15802
rect 1970 15750 1972 15802
rect 1996 15750 2034 15802
rect 2034 15750 2046 15802
rect 2046 15750 2052 15802
rect 2076 15750 2098 15802
rect 2098 15750 2110 15802
rect 2110 15750 2132 15802
rect 2156 15750 2162 15802
rect 2162 15750 2174 15802
rect 2174 15750 2212 15802
rect 2236 15750 2238 15802
rect 2238 15750 2290 15802
rect 2290 15750 2292 15802
rect 1916 15748 1972 15750
rect 1996 15748 2052 15750
rect 2076 15748 2132 15750
rect 2156 15748 2212 15750
rect 2236 15748 2292 15750
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 1916 14662 1918 14714
rect 1918 14662 1970 14714
rect 1970 14662 1972 14714
rect 1996 14662 2034 14714
rect 2034 14662 2046 14714
rect 2046 14662 2052 14714
rect 2076 14662 2098 14714
rect 2098 14662 2110 14714
rect 2110 14662 2132 14714
rect 2156 14662 2162 14714
rect 2162 14662 2174 14714
rect 2174 14662 2212 14714
rect 2236 14662 2238 14714
rect 2238 14662 2290 14714
rect 2290 14662 2292 14714
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 2656 15258 2712 15260
rect 2736 15258 2792 15260
rect 2816 15258 2872 15260
rect 2896 15258 2952 15260
rect 2976 15258 3032 15260
rect 2656 15206 2658 15258
rect 2658 15206 2710 15258
rect 2710 15206 2712 15258
rect 2736 15206 2774 15258
rect 2774 15206 2786 15258
rect 2786 15206 2792 15258
rect 2816 15206 2838 15258
rect 2838 15206 2850 15258
rect 2850 15206 2872 15258
rect 2896 15206 2902 15258
rect 2902 15206 2914 15258
rect 2914 15206 2952 15258
rect 2976 15206 2978 15258
rect 2978 15206 3030 15258
rect 3030 15206 3032 15258
rect 2656 15204 2712 15206
rect 2736 15204 2792 15206
rect 2816 15204 2872 15206
rect 2896 15204 2952 15206
rect 2976 15204 3032 15206
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 1916 13574 1918 13626
rect 1918 13574 1970 13626
rect 1970 13574 1972 13626
rect 1996 13574 2034 13626
rect 2034 13574 2046 13626
rect 2046 13574 2052 13626
rect 2076 13574 2098 13626
rect 2098 13574 2110 13626
rect 2110 13574 2132 13626
rect 2156 13574 2162 13626
rect 2162 13574 2174 13626
rect 2174 13574 2212 13626
rect 2236 13574 2238 13626
rect 2238 13574 2290 13626
rect 2290 13574 2292 13626
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 2656 14170 2712 14172
rect 2736 14170 2792 14172
rect 2816 14170 2872 14172
rect 2896 14170 2952 14172
rect 2976 14170 3032 14172
rect 2656 14118 2658 14170
rect 2658 14118 2710 14170
rect 2710 14118 2712 14170
rect 2736 14118 2774 14170
rect 2774 14118 2786 14170
rect 2786 14118 2792 14170
rect 2816 14118 2838 14170
rect 2838 14118 2850 14170
rect 2850 14118 2872 14170
rect 2896 14118 2902 14170
rect 2902 14118 2914 14170
rect 2914 14118 2952 14170
rect 2976 14118 2978 14170
rect 2978 14118 3030 14170
rect 3030 14118 3032 14170
rect 2656 14116 2712 14118
rect 2736 14116 2792 14118
rect 2816 14116 2872 14118
rect 2896 14116 2952 14118
rect 2976 14116 3032 14118
rect 2656 13082 2712 13084
rect 2736 13082 2792 13084
rect 2816 13082 2872 13084
rect 2896 13082 2952 13084
rect 2976 13082 3032 13084
rect 2656 13030 2658 13082
rect 2658 13030 2710 13082
rect 2710 13030 2712 13082
rect 2736 13030 2774 13082
rect 2774 13030 2786 13082
rect 2786 13030 2792 13082
rect 2816 13030 2838 13082
rect 2838 13030 2850 13082
rect 2850 13030 2872 13082
rect 2896 13030 2902 13082
rect 2902 13030 2914 13082
rect 2914 13030 2952 13082
rect 2976 13030 2978 13082
rect 2978 13030 3030 13082
rect 3030 13030 3032 13082
rect 2656 13028 2712 13030
rect 2736 13028 2792 13030
rect 2816 13028 2872 13030
rect 2896 13028 2952 13030
rect 2976 13028 3032 13030
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 1916 12486 1918 12538
rect 1918 12486 1970 12538
rect 1970 12486 1972 12538
rect 1996 12486 2034 12538
rect 2034 12486 2046 12538
rect 2046 12486 2052 12538
rect 2076 12486 2098 12538
rect 2098 12486 2110 12538
rect 2110 12486 2132 12538
rect 2156 12486 2162 12538
rect 2162 12486 2174 12538
rect 2174 12486 2212 12538
rect 2236 12486 2238 12538
rect 2238 12486 2290 12538
rect 2290 12486 2292 12538
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 2656 11994 2712 11996
rect 2736 11994 2792 11996
rect 2816 11994 2872 11996
rect 2896 11994 2952 11996
rect 2976 11994 3032 11996
rect 2656 11942 2658 11994
rect 2658 11942 2710 11994
rect 2710 11942 2712 11994
rect 2736 11942 2774 11994
rect 2774 11942 2786 11994
rect 2786 11942 2792 11994
rect 2816 11942 2838 11994
rect 2838 11942 2850 11994
rect 2850 11942 2872 11994
rect 2896 11942 2902 11994
rect 2902 11942 2914 11994
rect 2914 11942 2952 11994
rect 2976 11942 2978 11994
rect 2978 11942 3030 11994
rect 3030 11942 3032 11994
rect 2656 11940 2712 11942
rect 2736 11940 2792 11942
rect 2816 11940 2872 11942
rect 2896 11940 2952 11942
rect 2976 11940 3032 11942
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 1916 11398 1918 11450
rect 1918 11398 1970 11450
rect 1970 11398 1972 11450
rect 1996 11398 2034 11450
rect 2034 11398 2046 11450
rect 2046 11398 2052 11450
rect 2076 11398 2098 11450
rect 2098 11398 2110 11450
rect 2110 11398 2132 11450
rect 2156 11398 2162 11450
rect 2162 11398 2174 11450
rect 2174 11398 2212 11450
rect 2236 11398 2238 11450
rect 2238 11398 2290 11450
rect 2290 11398 2292 11450
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 1916 10310 1918 10362
rect 1918 10310 1970 10362
rect 1970 10310 1972 10362
rect 1996 10310 2034 10362
rect 2034 10310 2046 10362
rect 2046 10310 2052 10362
rect 2076 10310 2098 10362
rect 2098 10310 2110 10362
rect 2110 10310 2132 10362
rect 2156 10310 2162 10362
rect 2162 10310 2174 10362
rect 2174 10310 2212 10362
rect 2236 10310 2238 10362
rect 2238 10310 2290 10362
rect 2290 10310 2292 10362
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 2656 10906 2712 10908
rect 2736 10906 2792 10908
rect 2816 10906 2872 10908
rect 2896 10906 2952 10908
rect 2976 10906 3032 10908
rect 2656 10854 2658 10906
rect 2658 10854 2710 10906
rect 2710 10854 2712 10906
rect 2736 10854 2774 10906
rect 2774 10854 2786 10906
rect 2786 10854 2792 10906
rect 2816 10854 2838 10906
rect 2838 10854 2850 10906
rect 2850 10854 2872 10906
rect 2896 10854 2902 10906
rect 2902 10854 2914 10906
rect 2914 10854 2952 10906
rect 2976 10854 2978 10906
rect 2978 10854 3030 10906
rect 3030 10854 3032 10906
rect 2656 10852 2712 10854
rect 2736 10852 2792 10854
rect 2816 10852 2872 10854
rect 2896 10852 2952 10854
rect 2976 10852 3032 10854
rect 2656 9818 2712 9820
rect 2736 9818 2792 9820
rect 2816 9818 2872 9820
rect 2896 9818 2952 9820
rect 2976 9818 3032 9820
rect 2656 9766 2658 9818
rect 2658 9766 2710 9818
rect 2710 9766 2712 9818
rect 2736 9766 2774 9818
rect 2774 9766 2786 9818
rect 2786 9766 2792 9818
rect 2816 9766 2838 9818
rect 2838 9766 2850 9818
rect 2850 9766 2872 9818
rect 2896 9766 2902 9818
rect 2902 9766 2914 9818
rect 2914 9766 2952 9818
rect 2976 9766 2978 9818
rect 2978 9766 3030 9818
rect 3030 9766 3032 9818
rect 2656 9764 2712 9766
rect 2736 9764 2792 9766
rect 2816 9764 2872 9766
rect 2896 9764 2952 9766
rect 2976 9764 3032 9766
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 1916 9222 1918 9274
rect 1918 9222 1970 9274
rect 1970 9222 1972 9274
rect 1996 9222 2034 9274
rect 2034 9222 2046 9274
rect 2046 9222 2052 9274
rect 2076 9222 2098 9274
rect 2098 9222 2110 9274
rect 2110 9222 2132 9274
rect 2156 9222 2162 9274
rect 2162 9222 2174 9274
rect 2174 9222 2212 9274
rect 2236 9222 2238 9274
rect 2238 9222 2290 9274
rect 2290 9222 2292 9274
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 2656 8730 2712 8732
rect 2736 8730 2792 8732
rect 2816 8730 2872 8732
rect 2896 8730 2952 8732
rect 2976 8730 3032 8732
rect 2656 8678 2658 8730
rect 2658 8678 2710 8730
rect 2710 8678 2712 8730
rect 2736 8678 2774 8730
rect 2774 8678 2786 8730
rect 2786 8678 2792 8730
rect 2816 8678 2838 8730
rect 2838 8678 2850 8730
rect 2850 8678 2872 8730
rect 2896 8678 2902 8730
rect 2902 8678 2914 8730
rect 2914 8678 2952 8730
rect 2976 8678 2978 8730
rect 2978 8678 3030 8730
rect 3030 8678 3032 8730
rect 2656 8676 2712 8678
rect 2736 8676 2792 8678
rect 2816 8676 2872 8678
rect 2896 8676 2952 8678
rect 2976 8676 3032 8678
rect 7916 19066 7972 19068
rect 7996 19066 8052 19068
rect 8076 19066 8132 19068
rect 8156 19066 8212 19068
rect 8236 19066 8292 19068
rect 7916 19014 7918 19066
rect 7918 19014 7970 19066
rect 7970 19014 7972 19066
rect 7996 19014 8034 19066
rect 8034 19014 8046 19066
rect 8046 19014 8052 19066
rect 8076 19014 8098 19066
rect 8098 19014 8110 19066
rect 8110 19014 8132 19066
rect 8156 19014 8162 19066
rect 8162 19014 8174 19066
rect 8174 19014 8212 19066
rect 8236 19014 8238 19066
rect 8238 19014 8290 19066
rect 8290 19014 8292 19066
rect 7916 19012 7972 19014
rect 7996 19012 8052 19014
rect 8076 19012 8132 19014
rect 8156 19012 8212 19014
rect 8236 19012 8292 19014
rect 6366 14340 6422 14376
rect 6366 14320 6368 14340
rect 6368 14320 6420 14340
rect 6420 14320 6422 14340
rect 2656 7642 2712 7644
rect 2736 7642 2792 7644
rect 2816 7642 2872 7644
rect 2896 7642 2952 7644
rect 2976 7642 3032 7644
rect 2656 7590 2658 7642
rect 2658 7590 2710 7642
rect 2710 7590 2712 7642
rect 2736 7590 2774 7642
rect 2774 7590 2786 7642
rect 2786 7590 2792 7642
rect 2816 7590 2838 7642
rect 2838 7590 2850 7642
rect 2850 7590 2872 7642
rect 2896 7590 2902 7642
rect 2902 7590 2914 7642
rect 2914 7590 2952 7642
rect 2976 7590 2978 7642
rect 2978 7590 3030 7642
rect 3030 7590 3032 7642
rect 2656 7588 2712 7590
rect 2736 7588 2792 7590
rect 2816 7588 2872 7590
rect 2896 7588 2952 7590
rect 2976 7588 3032 7590
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 2656 6554 2712 6556
rect 2736 6554 2792 6556
rect 2816 6554 2872 6556
rect 2896 6554 2952 6556
rect 2976 6554 3032 6556
rect 2656 6502 2658 6554
rect 2658 6502 2710 6554
rect 2710 6502 2712 6554
rect 2736 6502 2774 6554
rect 2774 6502 2786 6554
rect 2786 6502 2792 6554
rect 2816 6502 2838 6554
rect 2838 6502 2850 6554
rect 2850 6502 2872 6554
rect 2896 6502 2902 6554
rect 2902 6502 2914 6554
rect 2914 6502 2952 6554
rect 2976 6502 2978 6554
rect 2978 6502 3030 6554
rect 3030 6502 3032 6554
rect 2656 6500 2712 6502
rect 2736 6500 2792 6502
rect 2816 6500 2872 6502
rect 2896 6500 2952 6502
rect 2976 6500 3032 6502
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 1306 5208 1362 5264
rect 2656 5466 2712 5468
rect 2736 5466 2792 5468
rect 2816 5466 2872 5468
rect 2896 5466 2952 5468
rect 2976 5466 3032 5468
rect 2656 5414 2658 5466
rect 2658 5414 2710 5466
rect 2710 5414 2712 5466
rect 2736 5414 2774 5466
rect 2774 5414 2786 5466
rect 2786 5414 2792 5466
rect 2816 5414 2838 5466
rect 2838 5414 2850 5466
rect 2850 5414 2872 5466
rect 2896 5414 2902 5466
rect 2902 5414 2914 5466
rect 2914 5414 2952 5466
rect 2976 5414 2978 5466
rect 2978 5414 3030 5466
rect 3030 5414 3032 5466
rect 2656 5412 2712 5414
rect 2736 5412 2792 5414
rect 2816 5412 2872 5414
rect 2896 5412 2952 5414
rect 2976 5412 3032 5414
rect 5998 8472 6054 8528
rect 8656 18522 8712 18524
rect 8736 18522 8792 18524
rect 8816 18522 8872 18524
rect 8896 18522 8952 18524
rect 8976 18522 9032 18524
rect 8656 18470 8658 18522
rect 8658 18470 8710 18522
rect 8710 18470 8712 18522
rect 8736 18470 8774 18522
rect 8774 18470 8786 18522
rect 8786 18470 8792 18522
rect 8816 18470 8838 18522
rect 8838 18470 8850 18522
rect 8850 18470 8872 18522
rect 8896 18470 8902 18522
rect 8902 18470 8914 18522
rect 8914 18470 8952 18522
rect 8976 18470 8978 18522
rect 8978 18470 9030 18522
rect 9030 18470 9032 18522
rect 8656 18468 8712 18470
rect 8736 18468 8792 18470
rect 8816 18468 8872 18470
rect 8896 18468 8952 18470
rect 8976 18468 9032 18470
rect 7916 17978 7972 17980
rect 7996 17978 8052 17980
rect 8076 17978 8132 17980
rect 8156 17978 8212 17980
rect 8236 17978 8292 17980
rect 7916 17926 7918 17978
rect 7918 17926 7970 17978
rect 7970 17926 7972 17978
rect 7996 17926 8034 17978
rect 8034 17926 8046 17978
rect 8046 17926 8052 17978
rect 8076 17926 8098 17978
rect 8098 17926 8110 17978
rect 8110 17926 8132 17978
rect 8156 17926 8162 17978
rect 8162 17926 8174 17978
rect 8174 17926 8212 17978
rect 8236 17926 8238 17978
rect 8238 17926 8290 17978
rect 8290 17926 8292 17978
rect 7916 17924 7972 17926
rect 7996 17924 8052 17926
rect 8076 17924 8132 17926
rect 8156 17924 8212 17926
rect 8236 17924 8292 17926
rect 8656 17434 8712 17436
rect 8736 17434 8792 17436
rect 8816 17434 8872 17436
rect 8896 17434 8952 17436
rect 8976 17434 9032 17436
rect 8656 17382 8658 17434
rect 8658 17382 8710 17434
rect 8710 17382 8712 17434
rect 8736 17382 8774 17434
rect 8774 17382 8786 17434
rect 8786 17382 8792 17434
rect 8816 17382 8838 17434
rect 8838 17382 8850 17434
rect 8850 17382 8872 17434
rect 8896 17382 8902 17434
rect 8902 17382 8914 17434
rect 8914 17382 8952 17434
rect 8976 17382 8978 17434
rect 8978 17382 9030 17434
rect 9030 17382 9032 17434
rect 8656 17380 8712 17382
rect 8736 17380 8792 17382
rect 8816 17380 8872 17382
rect 8896 17380 8952 17382
rect 8976 17380 9032 17382
rect 7916 16890 7972 16892
rect 7996 16890 8052 16892
rect 8076 16890 8132 16892
rect 8156 16890 8212 16892
rect 8236 16890 8292 16892
rect 7916 16838 7918 16890
rect 7918 16838 7970 16890
rect 7970 16838 7972 16890
rect 7996 16838 8034 16890
rect 8034 16838 8046 16890
rect 8046 16838 8052 16890
rect 8076 16838 8098 16890
rect 8098 16838 8110 16890
rect 8110 16838 8132 16890
rect 8156 16838 8162 16890
rect 8162 16838 8174 16890
rect 8174 16838 8212 16890
rect 8236 16838 8238 16890
rect 8238 16838 8290 16890
rect 8290 16838 8292 16890
rect 7916 16836 7972 16838
rect 7996 16836 8052 16838
rect 8076 16836 8132 16838
rect 8156 16836 8212 16838
rect 8236 16836 8292 16838
rect 8656 16346 8712 16348
rect 8736 16346 8792 16348
rect 8816 16346 8872 16348
rect 8896 16346 8952 16348
rect 8976 16346 9032 16348
rect 8656 16294 8658 16346
rect 8658 16294 8710 16346
rect 8710 16294 8712 16346
rect 8736 16294 8774 16346
rect 8774 16294 8786 16346
rect 8786 16294 8792 16346
rect 8816 16294 8838 16346
rect 8838 16294 8850 16346
rect 8850 16294 8872 16346
rect 8896 16294 8902 16346
rect 8902 16294 8914 16346
rect 8914 16294 8952 16346
rect 8976 16294 8978 16346
rect 8978 16294 9030 16346
rect 9030 16294 9032 16346
rect 8656 16292 8712 16294
rect 8736 16292 8792 16294
rect 8816 16292 8872 16294
rect 8896 16292 8952 16294
rect 8976 16292 9032 16294
rect 7916 15802 7972 15804
rect 7996 15802 8052 15804
rect 8076 15802 8132 15804
rect 8156 15802 8212 15804
rect 8236 15802 8292 15804
rect 7916 15750 7918 15802
rect 7918 15750 7970 15802
rect 7970 15750 7972 15802
rect 7996 15750 8034 15802
rect 8034 15750 8046 15802
rect 8046 15750 8052 15802
rect 8076 15750 8098 15802
rect 8098 15750 8110 15802
rect 8110 15750 8132 15802
rect 8156 15750 8162 15802
rect 8162 15750 8174 15802
rect 8174 15750 8212 15802
rect 8236 15750 8238 15802
rect 8238 15750 8290 15802
rect 8290 15750 8292 15802
rect 7916 15748 7972 15750
rect 7996 15748 8052 15750
rect 8076 15748 8132 15750
rect 8156 15748 8212 15750
rect 8236 15748 8292 15750
rect 7916 14714 7972 14716
rect 7996 14714 8052 14716
rect 8076 14714 8132 14716
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 7916 14662 7918 14714
rect 7918 14662 7970 14714
rect 7970 14662 7972 14714
rect 7996 14662 8034 14714
rect 8034 14662 8046 14714
rect 8046 14662 8052 14714
rect 8076 14662 8098 14714
rect 8098 14662 8110 14714
rect 8110 14662 8132 14714
rect 8156 14662 8162 14714
rect 8162 14662 8174 14714
rect 8174 14662 8212 14714
rect 8236 14662 8238 14714
rect 8238 14662 8290 14714
rect 8290 14662 8292 14714
rect 7916 14660 7972 14662
rect 7996 14660 8052 14662
rect 8076 14660 8132 14662
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 8656 15258 8712 15260
rect 8736 15258 8792 15260
rect 8816 15258 8872 15260
rect 8896 15258 8952 15260
rect 8976 15258 9032 15260
rect 8656 15206 8658 15258
rect 8658 15206 8710 15258
rect 8710 15206 8712 15258
rect 8736 15206 8774 15258
rect 8774 15206 8786 15258
rect 8786 15206 8792 15258
rect 8816 15206 8838 15258
rect 8838 15206 8850 15258
rect 8850 15206 8872 15258
rect 8896 15206 8902 15258
rect 8902 15206 8914 15258
rect 8914 15206 8952 15258
rect 8976 15206 8978 15258
rect 8978 15206 9030 15258
rect 9030 15206 9032 15258
rect 8656 15204 8712 15206
rect 8736 15204 8792 15206
rect 8816 15204 8872 15206
rect 8896 15204 8952 15206
rect 8976 15204 9032 15206
rect 8758 14340 8814 14376
rect 8758 14320 8760 14340
rect 8760 14320 8812 14340
rect 8812 14320 8814 14340
rect 8656 14170 8712 14172
rect 8736 14170 8792 14172
rect 8816 14170 8872 14172
rect 8896 14170 8952 14172
rect 8976 14170 9032 14172
rect 8656 14118 8658 14170
rect 8658 14118 8710 14170
rect 8710 14118 8712 14170
rect 8736 14118 8774 14170
rect 8774 14118 8786 14170
rect 8786 14118 8792 14170
rect 8816 14118 8838 14170
rect 8838 14118 8850 14170
rect 8850 14118 8872 14170
rect 8896 14118 8902 14170
rect 8902 14118 8914 14170
rect 8914 14118 8952 14170
rect 8976 14118 8978 14170
rect 8978 14118 9030 14170
rect 9030 14118 9032 14170
rect 8656 14116 8712 14118
rect 8736 14116 8792 14118
rect 8816 14116 8872 14118
rect 8896 14116 8952 14118
rect 8976 14116 9032 14118
rect 7916 13626 7972 13628
rect 7996 13626 8052 13628
rect 8076 13626 8132 13628
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 7916 13574 7918 13626
rect 7918 13574 7970 13626
rect 7970 13574 7972 13626
rect 7996 13574 8034 13626
rect 8034 13574 8046 13626
rect 8046 13574 8052 13626
rect 8076 13574 8098 13626
rect 8098 13574 8110 13626
rect 8110 13574 8132 13626
rect 8156 13574 8162 13626
rect 8162 13574 8174 13626
rect 8174 13574 8212 13626
rect 8236 13574 8238 13626
rect 8238 13574 8290 13626
rect 8290 13574 8292 13626
rect 7916 13572 7972 13574
rect 7996 13572 8052 13574
rect 8076 13572 8132 13574
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 8656 13082 8712 13084
rect 8736 13082 8792 13084
rect 8816 13082 8872 13084
rect 8896 13082 8952 13084
rect 8976 13082 9032 13084
rect 8656 13030 8658 13082
rect 8658 13030 8710 13082
rect 8710 13030 8712 13082
rect 8736 13030 8774 13082
rect 8774 13030 8786 13082
rect 8786 13030 8792 13082
rect 8816 13030 8838 13082
rect 8838 13030 8850 13082
rect 8850 13030 8872 13082
rect 8896 13030 8902 13082
rect 8902 13030 8914 13082
rect 8914 13030 8952 13082
rect 8976 13030 8978 13082
rect 8978 13030 9030 13082
rect 9030 13030 9032 13082
rect 8656 13028 8712 13030
rect 8736 13028 8792 13030
rect 8816 13028 8872 13030
rect 8896 13028 8952 13030
rect 8976 13028 9032 13030
rect 7916 12538 7972 12540
rect 7996 12538 8052 12540
rect 8076 12538 8132 12540
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 7916 12486 7918 12538
rect 7918 12486 7970 12538
rect 7970 12486 7972 12538
rect 7996 12486 8034 12538
rect 8034 12486 8046 12538
rect 8046 12486 8052 12538
rect 8076 12486 8098 12538
rect 8098 12486 8110 12538
rect 8110 12486 8132 12538
rect 8156 12486 8162 12538
rect 8162 12486 8174 12538
rect 8174 12486 8212 12538
rect 8236 12486 8238 12538
rect 8238 12486 8290 12538
rect 8290 12486 8292 12538
rect 7916 12484 7972 12486
rect 7996 12484 8052 12486
rect 8076 12484 8132 12486
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 7916 11450 7972 11452
rect 7996 11450 8052 11452
rect 8076 11450 8132 11452
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 7916 11398 7918 11450
rect 7918 11398 7970 11450
rect 7970 11398 7972 11450
rect 7996 11398 8034 11450
rect 8034 11398 8046 11450
rect 8046 11398 8052 11450
rect 8076 11398 8098 11450
rect 8098 11398 8110 11450
rect 8110 11398 8132 11450
rect 8156 11398 8162 11450
rect 8162 11398 8174 11450
rect 8174 11398 8212 11450
rect 8236 11398 8238 11450
rect 8238 11398 8290 11450
rect 8290 11398 8292 11450
rect 7916 11396 7972 11398
rect 7996 11396 8052 11398
rect 8076 11396 8132 11398
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 8656 11994 8712 11996
rect 8736 11994 8792 11996
rect 8816 11994 8872 11996
rect 8896 11994 8952 11996
rect 8976 11994 9032 11996
rect 8656 11942 8658 11994
rect 8658 11942 8710 11994
rect 8710 11942 8712 11994
rect 8736 11942 8774 11994
rect 8774 11942 8786 11994
rect 8786 11942 8792 11994
rect 8816 11942 8838 11994
rect 8838 11942 8850 11994
rect 8850 11942 8872 11994
rect 8896 11942 8902 11994
rect 8902 11942 8914 11994
rect 8914 11942 8952 11994
rect 8976 11942 8978 11994
rect 8978 11942 9030 11994
rect 9030 11942 9032 11994
rect 8656 11940 8712 11942
rect 8736 11940 8792 11942
rect 8816 11940 8872 11942
rect 8896 11940 8952 11942
rect 8976 11940 9032 11942
rect 7916 10362 7972 10364
rect 7996 10362 8052 10364
rect 8076 10362 8132 10364
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 7916 10310 7918 10362
rect 7918 10310 7970 10362
rect 7970 10310 7972 10362
rect 7996 10310 8034 10362
rect 8034 10310 8046 10362
rect 8046 10310 8052 10362
rect 8076 10310 8098 10362
rect 8098 10310 8110 10362
rect 8110 10310 8132 10362
rect 8156 10310 8162 10362
rect 8162 10310 8174 10362
rect 8174 10310 8212 10362
rect 8236 10310 8238 10362
rect 8238 10310 8290 10362
rect 8290 10310 8292 10362
rect 7916 10308 7972 10310
rect 7996 10308 8052 10310
rect 8076 10308 8132 10310
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 8656 10906 8712 10908
rect 8736 10906 8792 10908
rect 8816 10906 8872 10908
rect 8896 10906 8952 10908
rect 8976 10906 9032 10908
rect 8656 10854 8658 10906
rect 8658 10854 8710 10906
rect 8710 10854 8712 10906
rect 8736 10854 8774 10906
rect 8774 10854 8786 10906
rect 8786 10854 8792 10906
rect 8816 10854 8838 10906
rect 8838 10854 8850 10906
rect 8850 10854 8872 10906
rect 8896 10854 8902 10906
rect 8902 10854 8914 10906
rect 8914 10854 8952 10906
rect 8976 10854 8978 10906
rect 8978 10854 9030 10906
rect 9030 10854 9032 10906
rect 8656 10852 8712 10854
rect 8736 10852 8792 10854
rect 8816 10852 8872 10854
rect 8896 10852 8952 10854
rect 8976 10852 9032 10854
rect 8656 9818 8712 9820
rect 8736 9818 8792 9820
rect 8816 9818 8872 9820
rect 8896 9818 8952 9820
rect 8976 9818 9032 9820
rect 8656 9766 8658 9818
rect 8658 9766 8710 9818
rect 8710 9766 8712 9818
rect 8736 9766 8774 9818
rect 8774 9766 8786 9818
rect 8786 9766 8792 9818
rect 8816 9766 8838 9818
rect 8838 9766 8850 9818
rect 8850 9766 8872 9818
rect 8896 9766 8902 9818
rect 8902 9766 8914 9818
rect 8914 9766 8952 9818
rect 8976 9766 8978 9818
rect 8978 9766 9030 9818
rect 9030 9766 9032 9818
rect 8656 9764 8712 9766
rect 8736 9764 8792 9766
rect 8816 9764 8872 9766
rect 8896 9764 8952 9766
rect 8976 9764 9032 9766
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 8076 9274 8132 9276
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 7916 9222 7918 9274
rect 7918 9222 7970 9274
rect 7970 9222 7972 9274
rect 7996 9222 8034 9274
rect 8034 9222 8046 9274
rect 8046 9222 8052 9274
rect 8076 9222 8098 9274
rect 8098 9222 8110 9274
rect 8110 9222 8132 9274
rect 8156 9222 8162 9274
rect 8162 9222 8174 9274
rect 8174 9222 8212 9274
rect 8236 9222 8238 9274
rect 8238 9222 8290 9274
rect 8290 9222 8292 9274
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 8076 9220 8132 9222
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 8656 8730 8712 8732
rect 8736 8730 8792 8732
rect 8816 8730 8872 8732
rect 8896 8730 8952 8732
rect 8976 8730 9032 8732
rect 8656 8678 8658 8730
rect 8658 8678 8710 8730
rect 8710 8678 8712 8730
rect 8736 8678 8774 8730
rect 8774 8678 8786 8730
rect 8786 8678 8792 8730
rect 8816 8678 8838 8730
rect 8838 8678 8850 8730
rect 8850 8678 8872 8730
rect 8896 8678 8902 8730
rect 8902 8678 8914 8730
rect 8914 8678 8952 8730
rect 8976 8678 8978 8730
rect 8978 8678 9030 8730
rect 9030 8678 9032 8730
rect 8656 8676 8712 8678
rect 8736 8676 8792 8678
rect 8816 8676 8872 8678
rect 8896 8676 8952 8678
rect 8976 8676 9032 8678
rect 8758 8472 8814 8528
rect 8656 7642 8712 7644
rect 8736 7642 8792 7644
rect 8816 7642 8872 7644
rect 8896 7642 8952 7644
rect 8976 7642 9032 7644
rect 8656 7590 8658 7642
rect 8658 7590 8710 7642
rect 8710 7590 8712 7642
rect 8736 7590 8774 7642
rect 8774 7590 8786 7642
rect 8786 7590 8792 7642
rect 8816 7590 8838 7642
rect 8838 7590 8850 7642
rect 8850 7590 8872 7642
rect 8896 7590 8902 7642
rect 8902 7590 8914 7642
rect 8914 7590 8952 7642
rect 8976 7590 8978 7642
rect 8978 7590 9030 7642
rect 9030 7590 9032 7642
rect 8656 7588 8712 7590
rect 8736 7588 8792 7590
rect 8816 7588 8872 7590
rect 8896 7588 8952 7590
rect 8976 7588 9032 7590
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 10046 14320 10102 14376
rect 9862 8472 9918 8528
rect 8656 6554 8712 6556
rect 8736 6554 8792 6556
rect 8816 6554 8872 6556
rect 8896 6554 8952 6556
rect 8976 6554 9032 6556
rect 8656 6502 8658 6554
rect 8658 6502 8710 6554
rect 8710 6502 8712 6554
rect 8736 6502 8774 6554
rect 8774 6502 8786 6554
rect 8786 6502 8792 6554
rect 8816 6502 8838 6554
rect 8838 6502 8850 6554
rect 8850 6502 8872 6554
rect 8896 6502 8902 6554
rect 8902 6502 8914 6554
rect 8914 6502 8952 6554
rect 8976 6502 8978 6554
rect 8978 6502 9030 6554
rect 9030 6502 9032 6554
rect 8656 6500 8712 6502
rect 8736 6500 8792 6502
rect 8816 6500 8872 6502
rect 8896 6500 8952 6502
rect 8976 6500 9032 6502
rect 11334 11056 11390 11112
rect 8656 5466 8712 5468
rect 8736 5466 8792 5468
rect 8816 5466 8872 5468
rect 8896 5466 8952 5468
rect 8976 5466 9032 5468
rect 8656 5414 8658 5466
rect 8658 5414 8710 5466
rect 8710 5414 8712 5466
rect 8736 5414 8774 5466
rect 8774 5414 8786 5466
rect 8786 5414 8792 5466
rect 8816 5414 8838 5466
rect 8838 5414 8850 5466
rect 8850 5414 8872 5466
rect 8896 5414 8902 5466
rect 8902 5414 8914 5466
rect 8914 5414 8952 5466
rect 8976 5414 8978 5466
rect 8978 5414 9030 5466
rect 9030 5414 9032 5466
rect 8656 5412 8712 5414
rect 8736 5412 8792 5414
rect 8816 5412 8872 5414
rect 8896 5412 8952 5414
rect 8976 5412 9032 5414
rect 13916 19066 13972 19068
rect 13996 19066 14052 19068
rect 14076 19066 14132 19068
rect 14156 19066 14212 19068
rect 14236 19066 14292 19068
rect 13916 19014 13918 19066
rect 13918 19014 13970 19066
rect 13970 19014 13972 19066
rect 13996 19014 14034 19066
rect 14034 19014 14046 19066
rect 14046 19014 14052 19066
rect 14076 19014 14098 19066
rect 14098 19014 14110 19066
rect 14110 19014 14132 19066
rect 14156 19014 14162 19066
rect 14162 19014 14174 19066
rect 14174 19014 14212 19066
rect 14236 19014 14238 19066
rect 14238 19014 14290 19066
rect 14290 19014 14292 19066
rect 13916 19012 13972 19014
rect 13996 19012 14052 19014
rect 14076 19012 14132 19014
rect 14156 19012 14212 19014
rect 14236 19012 14292 19014
rect 14656 18522 14712 18524
rect 14736 18522 14792 18524
rect 14816 18522 14872 18524
rect 14896 18522 14952 18524
rect 14976 18522 15032 18524
rect 14656 18470 14658 18522
rect 14658 18470 14710 18522
rect 14710 18470 14712 18522
rect 14736 18470 14774 18522
rect 14774 18470 14786 18522
rect 14786 18470 14792 18522
rect 14816 18470 14838 18522
rect 14838 18470 14850 18522
rect 14850 18470 14872 18522
rect 14896 18470 14902 18522
rect 14902 18470 14914 18522
rect 14914 18470 14952 18522
rect 14976 18470 14978 18522
rect 14978 18470 15030 18522
rect 15030 18470 15032 18522
rect 14656 18468 14712 18470
rect 14736 18468 14792 18470
rect 14816 18468 14872 18470
rect 14896 18468 14952 18470
rect 14976 18468 15032 18470
rect 13916 17978 13972 17980
rect 13996 17978 14052 17980
rect 14076 17978 14132 17980
rect 14156 17978 14212 17980
rect 14236 17978 14292 17980
rect 13916 17926 13918 17978
rect 13918 17926 13970 17978
rect 13970 17926 13972 17978
rect 13996 17926 14034 17978
rect 14034 17926 14046 17978
rect 14046 17926 14052 17978
rect 14076 17926 14098 17978
rect 14098 17926 14110 17978
rect 14110 17926 14132 17978
rect 14156 17926 14162 17978
rect 14162 17926 14174 17978
rect 14174 17926 14212 17978
rect 14236 17926 14238 17978
rect 14238 17926 14290 17978
rect 14290 17926 14292 17978
rect 13916 17924 13972 17926
rect 13996 17924 14052 17926
rect 14076 17924 14132 17926
rect 14156 17924 14212 17926
rect 14236 17924 14292 17926
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 14156 16890 14212 16892
rect 14236 16890 14292 16892
rect 13916 16838 13918 16890
rect 13918 16838 13970 16890
rect 13970 16838 13972 16890
rect 13996 16838 14034 16890
rect 14034 16838 14046 16890
rect 14046 16838 14052 16890
rect 14076 16838 14098 16890
rect 14098 16838 14110 16890
rect 14110 16838 14132 16890
rect 14156 16838 14162 16890
rect 14162 16838 14174 16890
rect 14174 16838 14212 16890
rect 14236 16838 14238 16890
rect 14238 16838 14290 16890
rect 14290 16838 14292 16890
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 14156 16836 14212 16838
rect 14236 16836 14292 16838
rect 14656 17434 14712 17436
rect 14736 17434 14792 17436
rect 14816 17434 14872 17436
rect 14896 17434 14952 17436
rect 14976 17434 15032 17436
rect 14656 17382 14658 17434
rect 14658 17382 14710 17434
rect 14710 17382 14712 17434
rect 14736 17382 14774 17434
rect 14774 17382 14786 17434
rect 14786 17382 14792 17434
rect 14816 17382 14838 17434
rect 14838 17382 14850 17434
rect 14850 17382 14872 17434
rect 14896 17382 14902 17434
rect 14902 17382 14914 17434
rect 14914 17382 14952 17434
rect 14976 17382 14978 17434
rect 14978 17382 15030 17434
rect 15030 17382 15032 17434
rect 14656 17380 14712 17382
rect 14736 17380 14792 17382
rect 14816 17380 14872 17382
rect 14896 17380 14952 17382
rect 14976 17380 15032 17382
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 14156 15802 14212 15804
rect 14236 15802 14292 15804
rect 13916 15750 13918 15802
rect 13918 15750 13970 15802
rect 13970 15750 13972 15802
rect 13996 15750 14034 15802
rect 14034 15750 14046 15802
rect 14046 15750 14052 15802
rect 14076 15750 14098 15802
rect 14098 15750 14110 15802
rect 14110 15750 14132 15802
rect 14156 15750 14162 15802
rect 14162 15750 14174 15802
rect 14174 15750 14212 15802
rect 14236 15750 14238 15802
rect 14238 15750 14290 15802
rect 14290 15750 14292 15802
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 14156 15748 14212 15750
rect 14236 15748 14292 15750
rect 14656 16346 14712 16348
rect 14736 16346 14792 16348
rect 14816 16346 14872 16348
rect 14896 16346 14952 16348
rect 14976 16346 15032 16348
rect 14656 16294 14658 16346
rect 14658 16294 14710 16346
rect 14710 16294 14712 16346
rect 14736 16294 14774 16346
rect 14774 16294 14786 16346
rect 14786 16294 14792 16346
rect 14816 16294 14838 16346
rect 14838 16294 14850 16346
rect 14850 16294 14872 16346
rect 14896 16294 14902 16346
rect 14902 16294 14914 16346
rect 14914 16294 14952 16346
rect 14976 16294 14978 16346
rect 14978 16294 15030 16346
rect 15030 16294 15032 16346
rect 14656 16292 14712 16294
rect 14736 16292 14792 16294
rect 14816 16292 14872 16294
rect 14896 16292 14952 16294
rect 14976 16292 15032 16294
rect 13542 14340 13598 14376
rect 13542 14320 13544 14340
rect 13544 14320 13596 14340
rect 13596 14320 13598 14340
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 14156 14714 14212 14716
rect 14236 14714 14292 14716
rect 13916 14662 13918 14714
rect 13918 14662 13970 14714
rect 13970 14662 13972 14714
rect 13996 14662 14034 14714
rect 14034 14662 14046 14714
rect 14046 14662 14052 14714
rect 14076 14662 14098 14714
rect 14098 14662 14110 14714
rect 14110 14662 14132 14714
rect 14156 14662 14162 14714
rect 14162 14662 14174 14714
rect 14174 14662 14212 14714
rect 14236 14662 14238 14714
rect 14238 14662 14290 14714
rect 14290 14662 14292 14714
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 14156 14660 14212 14662
rect 14236 14660 14292 14662
rect 14656 15258 14712 15260
rect 14736 15258 14792 15260
rect 14816 15258 14872 15260
rect 14896 15258 14952 15260
rect 14976 15258 15032 15260
rect 14656 15206 14658 15258
rect 14658 15206 14710 15258
rect 14710 15206 14712 15258
rect 14736 15206 14774 15258
rect 14774 15206 14786 15258
rect 14786 15206 14792 15258
rect 14816 15206 14838 15258
rect 14838 15206 14850 15258
rect 14850 15206 14872 15258
rect 14896 15206 14902 15258
rect 14902 15206 14914 15258
rect 14914 15206 14952 15258
rect 14976 15206 14978 15258
rect 14978 15206 15030 15258
rect 15030 15206 15032 15258
rect 14656 15204 14712 15206
rect 14736 15204 14792 15206
rect 14816 15204 14872 15206
rect 14896 15204 14952 15206
rect 14976 15204 15032 15206
rect 14656 14170 14712 14172
rect 14736 14170 14792 14172
rect 14816 14170 14872 14172
rect 14896 14170 14952 14172
rect 14976 14170 15032 14172
rect 14656 14118 14658 14170
rect 14658 14118 14710 14170
rect 14710 14118 14712 14170
rect 14736 14118 14774 14170
rect 14774 14118 14786 14170
rect 14786 14118 14792 14170
rect 14816 14118 14838 14170
rect 14838 14118 14850 14170
rect 14850 14118 14872 14170
rect 14896 14118 14902 14170
rect 14902 14118 14914 14170
rect 14914 14118 14952 14170
rect 14976 14118 14978 14170
rect 14978 14118 15030 14170
rect 15030 14118 15032 14170
rect 14656 14116 14712 14118
rect 14736 14116 14792 14118
rect 14816 14116 14872 14118
rect 14896 14116 14952 14118
rect 14976 14116 15032 14118
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 14156 13626 14212 13628
rect 14236 13626 14292 13628
rect 13916 13574 13918 13626
rect 13918 13574 13970 13626
rect 13970 13574 13972 13626
rect 13996 13574 14034 13626
rect 14034 13574 14046 13626
rect 14046 13574 14052 13626
rect 14076 13574 14098 13626
rect 14098 13574 14110 13626
rect 14110 13574 14132 13626
rect 14156 13574 14162 13626
rect 14162 13574 14174 13626
rect 14174 13574 14212 13626
rect 14236 13574 14238 13626
rect 14238 13574 14290 13626
rect 14290 13574 14292 13626
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 14156 13572 14212 13574
rect 14236 13572 14292 13574
rect 14656 13082 14712 13084
rect 14736 13082 14792 13084
rect 14816 13082 14872 13084
rect 14896 13082 14952 13084
rect 14976 13082 15032 13084
rect 14656 13030 14658 13082
rect 14658 13030 14710 13082
rect 14710 13030 14712 13082
rect 14736 13030 14774 13082
rect 14774 13030 14786 13082
rect 14786 13030 14792 13082
rect 14816 13030 14838 13082
rect 14838 13030 14850 13082
rect 14850 13030 14872 13082
rect 14896 13030 14902 13082
rect 14902 13030 14914 13082
rect 14914 13030 14952 13082
rect 14976 13030 14978 13082
rect 14978 13030 15030 13082
rect 15030 13030 15032 13082
rect 14656 13028 14712 13030
rect 14736 13028 14792 13030
rect 14816 13028 14872 13030
rect 14896 13028 14952 13030
rect 14976 13028 15032 13030
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 14156 12538 14212 12540
rect 14236 12538 14292 12540
rect 13916 12486 13918 12538
rect 13918 12486 13970 12538
rect 13970 12486 13972 12538
rect 13996 12486 14034 12538
rect 14034 12486 14046 12538
rect 14046 12486 14052 12538
rect 14076 12486 14098 12538
rect 14098 12486 14110 12538
rect 14110 12486 14132 12538
rect 14156 12486 14162 12538
rect 14162 12486 14174 12538
rect 14174 12486 14212 12538
rect 14236 12486 14238 12538
rect 14238 12486 14290 12538
rect 14290 12486 14292 12538
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 14156 12484 14212 12486
rect 14236 12484 14292 12486
rect 14656 11994 14712 11996
rect 14736 11994 14792 11996
rect 14816 11994 14872 11996
rect 14896 11994 14952 11996
rect 14976 11994 15032 11996
rect 14656 11942 14658 11994
rect 14658 11942 14710 11994
rect 14710 11942 14712 11994
rect 14736 11942 14774 11994
rect 14774 11942 14786 11994
rect 14786 11942 14792 11994
rect 14816 11942 14838 11994
rect 14838 11942 14850 11994
rect 14850 11942 14872 11994
rect 14896 11942 14902 11994
rect 14902 11942 14914 11994
rect 14914 11942 14952 11994
rect 14976 11942 14978 11994
rect 14978 11942 15030 11994
rect 15030 11942 15032 11994
rect 14656 11940 14712 11942
rect 14736 11940 14792 11942
rect 14816 11940 14872 11942
rect 14896 11940 14952 11942
rect 14976 11940 15032 11942
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 14156 11450 14212 11452
rect 14236 11450 14292 11452
rect 13916 11398 13918 11450
rect 13918 11398 13970 11450
rect 13970 11398 13972 11450
rect 13996 11398 14034 11450
rect 14034 11398 14046 11450
rect 14046 11398 14052 11450
rect 14076 11398 14098 11450
rect 14098 11398 14110 11450
rect 14110 11398 14132 11450
rect 14156 11398 14162 11450
rect 14162 11398 14174 11450
rect 14174 11398 14212 11450
rect 14236 11398 14238 11450
rect 14238 11398 14290 11450
rect 14290 11398 14292 11450
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 14156 11396 14212 11398
rect 14236 11396 14292 11398
rect 14656 10906 14712 10908
rect 14736 10906 14792 10908
rect 14816 10906 14872 10908
rect 14896 10906 14952 10908
rect 14976 10906 15032 10908
rect 14656 10854 14658 10906
rect 14658 10854 14710 10906
rect 14710 10854 14712 10906
rect 14736 10854 14774 10906
rect 14774 10854 14786 10906
rect 14786 10854 14792 10906
rect 14816 10854 14838 10906
rect 14838 10854 14850 10906
rect 14850 10854 14872 10906
rect 14896 10854 14902 10906
rect 14902 10854 14914 10906
rect 14914 10854 14952 10906
rect 14976 10854 14978 10906
rect 14978 10854 15030 10906
rect 15030 10854 15032 10906
rect 14656 10852 14712 10854
rect 14736 10852 14792 10854
rect 14816 10852 14872 10854
rect 14896 10852 14952 10854
rect 14976 10852 15032 10854
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 14156 10362 14212 10364
rect 14236 10362 14292 10364
rect 13916 10310 13918 10362
rect 13918 10310 13970 10362
rect 13970 10310 13972 10362
rect 13996 10310 14034 10362
rect 14034 10310 14046 10362
rect 14046 10310 14052 10362
rect 14076 10310 14098 10362
rect 14098 10310 14110 10362
rect 14110 10310 14132 10362
rect 14156 10310 14162 10362
rect 14162 10310 14174 10362
rect 14174 10310 14212 10362
rect 14236 10310 14238 10362
rect 14238 10310 14290 10362
rect 14290 10310 14292 10362
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 14156 10308 14212 10310
rect 14236 10308 14292 10310
rect 14656 9818 14712 9820
rect 14736 9818 14792 9820
rect 14816 9818 14872 9820
rect 14896 9818 14952 9820
rect 14976 9818 15032 9820
rect 14656 9766 14658 9818
rect 14658 9766 14710 9818
rect 14710 9766 14712 9818
rect 14736 9766 14774 9818
rect 14774 9766 14786 9818
rect 14786 9766 14792 9818
rect 14816 9766 14838 9818
rect 14838 9766 14850 9818
rect 14850 9766 14872 9818
rect 14896 9766 14902 9818
rect 14902 9766 14914 9818
rect 14914 9766 14952 9818
rect 14976 9766 14978 9818
rect 14978 9766 15030 9818
rect 15030 9766 15032 9818
rect 14656 9764 14712 9766
rect 14736 9764 14792 9766
rect 14816 9764 14872 9766
rect 14896 9764 14952 9766
rect 14976 9764 15032 9766
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 14156 9274 14212 9276
rect 14236 9274 14292 9276
rect 13916 9222 13918 9274
rect 13918 9222 13970 9274
rect 13970 9222 13972 9274
rect 13996 9222 14034 9274
rect 14034 9222 14046 9274
rect 14046 9222 14052 9274
rect 14076 9222 14098 9274
rect 14098 9222 14110 9274
rect 14110 9222 14132 9274
rect 14156 9222 14162 9274
rect 14162 9222 14174 9274
rect 14174 9222 14212 9274
rect 14236 9222 14238 9274
rect 14238 9222 14290 9274
rect 14290 9222 14292 9274
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 14156 9220 14212 9222
rect 14236 9220 14292 9222
rect 13818 8472 13874 8528
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 14156 8186 14212 8188
rect 14236 8186 14292 8188
rect 13916 8134 13918 8186
rect 13918 8134 13970 8186
rect 13970 8134 13972 8186
rect 13996 8134 14034 8186
rect 14034 8134 14046 8186
rect 14046 8134 14052 8186
rect 14076 8134 14098 8186
rect 14098 8134 14110 8186
rect 14110 8134 14132 8186
rect 14156 8134 14162 8186
rect 14162 8134 14174 8186
rect 14174 8134 14212 8186
rect 14236 8134 14238 8186
rect 14238 8134 14290 8186
rect 14290 8134 14292 8186
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 14156 8132 14212 8134
rect 14236 8132 14292 8134
rect 14656 8730 14712 8732
rect 14736 8730 14792 8732
rect 14816 8730 14872 8732
rect 14896 8730 14952 8732
rect 14976 8730 15032 8732
rect 14656 8678 14658 8730
rect 14658 8678 14710 8730
rect 14710 8678 14712 8730
rect 14736 8678 14774 8730
rect 14774 8678 14786 8730
rect 14786 8678 14792 8730
rect 14816 8678 14838 8730
rect 14838 8678 14850 8730
rect 14850 8678 14872 8730
rect 14896 8678 14902 8730
rect 14902 8678 14914 8730
rect 14914 8678 14952 8730
rect 14976 8678 14978 8730
rect 14978 8678 15030 8730
rect 15030 8678 15032 8730
rect 14656 8676 14712 8678
rect 14736 8676 14792 8678
rect 14816 8676 14872 8678
rect 14896 8676 14952 8678
rect 14976 8676 15032 8678
rect 14646 8492 14702 8528
rect 14646 8472 14648 8492
rect 14648 8472 14700 8492
rect 14700 8472 14702 8492
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 14156 7098 14212 7100
rect 14236 7098 14292 7100
rect 13916 7046 13918 7098
rect 13918 7046 13970 7098
rect 13970 7046 13972 7098
rect 13996 7046 14034 7098
rect 14034 7046 14046 7098
rect 14046 7046 14052 7098
rect 14076 7046 14098 7098
rect 14098 7046 14110 7098
rect 14110 7046 14132 7098
rect 14156 7046 14162 7098
rect 14162 7046 14174 7098
rect 14174 7046 14212 7098
rect 14236 7046 14238 7098
rect 14238 7046 14290 7098
rect 14290 7046 14292 7098
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 14156 7044 14212 7046
rect 14236 7044 14292 7046
rect 14656 7642 14712 7644
rect 14736 7642 14792 7644
rect 14816 7642 14872 7644
rect 14896 7642 14952 7644
rect 14976 7642 15032 7644
rect 14656 7590 14658 7642
rect 14658 7590 14710 7642
rect 14710 7590 14712 7642
rect 14736 7590 14774 7642
rect 14774 7590 14786 7642
rect 14786 7590 14792 7642
rect 14816 7590 14838 7642
rect 14838 7590 14850 7642
rect 14850 7590 14872 7642
rect 14896 7590 14902 7642
rect 14902 7590 14914 7642
rect 14914 7590 14952 7642
rect 14976 7590 14978 7642
rect 14978 7590 15030 7642
rect 15030 7590 15032 7642
rect 14656 7588 14712 7590
rect 14736 7588 14792 7590
rect 14816 7588 14872 7590
rect 14896 7588 14952 7590
rect 14976 7588 15032 7590
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 14156 6010 14212 6012
rect 14236 6010 14292 6012
rect 13916 5958 13918 6010
rect 13918 5958 13970 6010
rect 13970 5958 13972 6010
rect 13996 5958 14034 6010
rect 14034 5958 14046 6010
rect 14046 5958 14052 6010
rect 14076 5958 14098 6010
rect 14098 5958 14110 6010
rect 14110 5958 14132 6010
rect 14156 5958 14162 6010
rect 14162 5958 14174 6010
rect 14174 5958 14212 6010
rect 14236 5958 14238 6010
rect 14238 5958 14290 6010
rect 14290 5958 14292 6010
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 14156 5956 14212 5958
rect 14236 5956 14292 5958
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 14656 6554 14712 6556
rect 14736 6554 14792 6556
rect 14816 6554 14872 6556
rect 14896 6554 14952 6556
rect 14976 6554 15032 6556
rect 14656 6502 14658 6554
rect 14658 6502 14710 6554
rect 14710 6502 14712 6554
rect 14736 6502 14774 6554
rect 14774 6502 14786 6554
rect 14786 6502 14792 6554
rect 14816 6502 14838 6554
rect 14838 6502 14850 6554
rect 14850 6502 14872 6554
rect 14896 6502 14902 6554
rect 14902 6502 14914 6554
rect 14914 6502 14952 6554
rect 14976 6502 14978 6554
rect 14978 6502 15030 6554
rect 15030 6502 15032 6554
rect 14656 6500 14712 6502
rect 14736 6500 14792 6502
rect 14816 6500 14872 6502
rect 14896 6500 14952 6502
rect 14976 6500 15032 6502
rect 16670 17992 16726 18048
rect 14656 5466 14712 5468
rect 14736 5466 14792 5468
rect 14816 5466 14872 5468
rect 14896 5466 14952 5468
rect 14976 5466 15032 5468
rect 14656 5414 14658 5466
rect 14658 5414 14710 5466
rect 14710 5414 14712 5466
rect 14736 5414 14774 5466
rect 14774 5414 14786 5466
rect 14786 5414 14792 5466
rect 14816 5414 14838 5466
rect 14838 5414 14850 5466
rect 14850 5414 14872 5466
rect 14896 5414 14902 5466
rect 14902 5414 14914 5466
rect 14914 5414 14952 5466
rect 14976 5414 14978 5466
rect 14978 5414 15030 5466
rect 15030 5414 15032 5466
rect 14656 5412 14712 5414
rect 14736 5412 14792 5414
rect 14816 5412 14872 5414
rect 14896 5412 14952 5414
rect 14976 5412 15032 5414
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 14156 4922 14212 4924
rect 14236 4922 14292 4924
rect 13916 4870 13918 4922
rect 13918 4870 13970 4922
rect 13970 4870 13972 4922
rect 13996 4870 14034 4922
rect 14034 4870 14046 4922
rect 14046 4870 14052 4922
rect 14076 4870 14098 4922
rect 14098 4870 14110 4922
rect 14110 4870 14132 4922
rect 14156 4870 14162 4922
rect 14162 4870 14174 4922
rect 14174 4870 14212 4922
rect 14236 4870 14238 4922
rect 14238 4870 14290 4922
rect 14290 4870 14292 4922
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 14156 4868 14212 4870
rect 14236 4868 14292 4870
rect 16578 5752 16634 5808
rect 2656 4378 2712 4380
rect 2736 4378 2792 4380
rect 2816 4378 2872 4380
rect 2896 4378 2952 4380
rect 2976 4378 3032 4380
rect 2656 4326 2658 4378
rect 2658 4326 2710 4378
rect 2710 4326 2712 4378
rect 2736 4326 2774 4378
rect 2774 4326 2786 4378
rect 2786 4326 2792 4378
rect 2816 4326 2838 4378
rect 2838 4326 2850 4378
rect 2850 4326 2872 4378
rect 2896 4326 2902 4378
rect 2902 4326 2914 4378
rect 2914 4326 2952 4378
rect 2976 4326 2978 4378
rect 2978 4326 3030 4378
rect 3030 4326 3032 4378
rect 2656 4324 2712 4326
rect 2736 4324 2792 4326
rect 2816 4324 2872 4326
rect 2896 4324 2952 4326
rect 2976 4324 3032 4326
rect 8656 4378 8712 4380
rect 8736 4378 8792 4380
rect 8816 4378 8872 4380
rect 8896 4378 8952 4380
rect 8976 4378 9032 4380
rect 8656 4326 8658 4378
rect 8658 4326 8710 4378
rect 8710 4326 8712 4378
rect 8736 4326 8774 4378
rect 8774 4326 8786 4378
rect 8786 4326 8792 4378
rect 8816 4326 8838 4378
rect 8838 4326 8850 4378
rect 8850 4326 8872 4378
rect 8896 4326 8902 4378
rect 8902 4326 8914 4378
rect 8914 4326 8952 4378
rect 8976 4326 8978 4378
rect 8978 4326 9030 4378
rect 9030 4326 9032 4378
rect 8656 4324 8712 4326
rect 8736 4324 8792 4326
rect 8816 4324 8872 4326
rect 8896 4324 8952 4326
rect 8976 4324 9032 4326
rect 14656 4378 14712 4380
rect 14736 4378 14792 4380
rect 14816 4378 14872 4380
rect 14896 4378 14952 4380
rect 14976 4378 15032 4380
rect 14656 4326 14658 4378
rect 14658 4326 14710 4378
rect 14710 4326 14712 4378
rect 14736 4326 14774 4378
rect 14774 4326 14786 4378
rect 14786 4326 14792 4378
rect 14816 4326 14838 4378
rect 14838 4326 14850 4378
rect 14850 4326 14872 4378
rect 14896 4326 14902 4378
rect 14902 4326 14914 4378
rect 14914 4326 14952 4378
rect 14976 4326 14978 4378
rect 14978 4326 15030 4378
rect 15030 4326 15032 4378
rect 14656 4324 14712 4326
rect 14736 4324 14792 4326
rect 14816 4324 14872 4326
rect 14896 4324 14952 4326
rect 14976 4324 15032 4326
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 14156 3834 14212 3836
rect 14236 3834 14292 3836
rect 13916 3782 13918 3834
rect 13918 3782 13970 3834
rect 13970 3782 13972 3834
rect 13996 3782 14034 3834
rect 14034 3782 14046 3834
rect 14046 3782 14052 3834
rect 14076 3782 14098 3834
rect 14098 3782 14110 3834
rect 14110 3782 14132 3834
rect 14156 3782 14162 3834
rect 14162 3782 14174 3834
rect 14174 3782 14212 3834
rect 14236 3782 14238 3834
rect 14238 3782 14290 3834
rect 14290 3782 14292 3834
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 14156 3780 14212 3782
rect 14236 3780 14292 3782
rect 2656 3290 2712 3292
rect 2736 3290 2792 3292
rect 2816 3290 2872 3292
rect 2896 3290 2952 3292
rect 2976 3290 3032 3292
rect 2656 3238 2658 3290
rect 2658 3238 2710 3290
rect 2710 3238 2712 3290
rect 2736 3238 2774 3290
rect 2774 3238 2786 3290
rect 2786 3238 2792 3290
rect 2816 3238 2838 3290
rect 2838 3238 2850 3290
rect 2850 3238 2872 3290
rect 2896 3238 2902 3290
rect 2902 3238 2914 3290
rect 2914 3238 2952 3290
rect 2976 3238 2978 3290
rect 2978 3238 3030 3290
rect 3030 3238 3032 3290
rect 2656 3236 2712 3238
rect 2736 3236 2792 3238
rect 2816 3236 2872 3238
rect 2896 3236 2952 3238
rect 2976 3236 3032 3238
rect 8656 3290 8712 3292
rect 8736 3290 8792 3292
rect 8816 3290 8872 3292
rect 8896 3290 8952 3292
rect 8976 3290 9032 3292
rect 8656 3238 8658 3290
rect 8658 3238 8710 3290
rect 8710 3238 8712 3290
rect 8736 3238 8774 3290
rect 8774 3238 8786 3290
rect 8786 3238 8792 3290
rect 8816 3238 8838 3290
rect 8838 3238 8850 3290
rect 8850 3238 8872 3290
rect 8896 3238 8902 3290
rect 8902 3238 8914 3290
rect 8914 3238 8952 3290
rect 8976 3238 8978 3290
rect 8978 3238 9030 3290
rect 9030 3238 9032 3290
rect 8656 3236 8712 3238
rect 8736 3236 8792 3238
rect 8816 3236 8872 3238
rect 8896 3236 8952 3238
rect 8976 3236 9032 3238
rect 14656 3290 14712 3292
rect 14736 3290 14792 3292
rect 14816 3290 14872 3292
rect 14896 3290 14952 3292
rect 14976 3290 15032 3292
rect 14656 3238 14658 3290
rect 14658 3238 14710 3290
rect 14710 3238 14712 3290
rect 14736 3238 14774 3290
rect 14774 3238 14786 3290
rect 14786 3238 14792 3290
rect 14816 3238 14838 3290
rect 14838 3238 14850 3290
rect 14850 3238 14872 3290
rect 14896 3238 14902 3290
rect 14902 3238 14914 3290
rect 14914 3238 14952 3290
rect 14976 3238 14978 3290
rect 14978 3238 15030 3290
rect 15030 3238 15032 3290
rect 14656 3236 14712 3238
rect 14736 3236 14792 3238
rect 14816 3236 14872 3238
rect 14896 3236 14952 3238
rect 14976 3236 15032 3238
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 14156 2746 14212 2748
rect 14236 2746 14292 2748
rect 13916 2694 13918 2746
rect 13918 2694 13970 2746
rect 13970 2694 13972 2746
rect 13996 2694 14034 2746
rect 14034 2694 14046 2746
rect 14046 2694 14052 2746
rect 14076 2694 14098 2746
rect 14098 2694 14110 2746
rect 14110 2694 14132 2746
rect 14156 2694 14162 2746
rect 14162 2694 14174 2746
rect 14174 2694 14212 2746
rect 14236 2694 14238 2746
rect 14238 2694 14290 2746
rect 14290 2694 14292 2746
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 14156 2692 14212 2694
rect 14236 2692 14292 2694
rect 2656 2202 2712 2204
rect 2736 2202 2792 2204
rect 2816 2202 2872 2204
rect 2896 2202 2952 2204
rect 2976 2202 3032 2204
rect 2656 2150 2658 2202
rect 2658 2150 2710 2202
rect 2710 2150 2712 2202
rect 2736 2150 2774 2202
rect 2774 2150 2786 2202
rect 2786 2150 2792 2202
rect 2816 2150 2838 2202
rect 2838 2150 2850 2202
rect 2850 2150 2872 2202
rect 2896 2150 2902 2202
rect 2902 2150 2914 2202
rect 2914 2150 2952 2202
rect 2976 2150 2978 2202
rect 2978 2150 3030 2202
rect 3030 2150 3032 2202
rect 2656 2148 2712 2150
rect 2736 2148 2792 2150
rect 2816 2148 2872 2150
rect 2896 2148 2952 2150
rect 2976 2148 3032 2150
rect 8656 2202 8712 2204
rect 8736 2202 8792 2204
rect 8816 2202 8872 2204
rect 8896 2202 8952 2204
rect 8976 2202 9032 2204
rect 8656 2150 8658 2202
rect 8658 2150 8710 2202
rect 8710 2150 8712 2202
rect 8736 2150 8774 2202
rect 8774 2150 8786 2202
rect 8786 2150 8792 2202
rect 8816 2150 8838 2202
rect 8838 2150 8850 2202
rect 8850 2150 8872 2202
rect 8896 2150 8902 2202
rect 8902 2150 8914 2202
rect 8914 2150 8952 2202
rect 8976 2150 8978 2202
rect 8978 2150 9030 2202
rect 9030 2150 9032 2202
rect 8656 2148 8712 2150
rect 8736 2148 8792 2150
rect 8816 2148 8872 2150
rect 8896 2148 8952 2150
rect 8976 2148 9032 2150
rect 14656 2202 14712 2204
rect 14736 2202 14792 2204
rect 14816 2202 14872 2204
rect 14896 2202 14952 2204
rect 14976 2202 15032 2204
rect 14656 2150 14658 2202
rect 14658 2150 14710 2202
rect 14710 2150 14712 2202
rect 14736 2150 14774 2202
rect 14774 2150 14786 2202
rect 14786 2150 14792 2202
rect 14816 2150 14838 2202
rect 14838 2150 14850 2202
rect 14850 2150 14872 2202
rect 14896 2150 14902 2202
rect 14902 2150 14914 2202
rect 14914 2150 14952 2202
rect 14976 2150 14978 2202
rect 14978 2150 15030 2202
rect 15030 2150 15032 2202
rect 14656 2148 14712 2150
rect 14736 2148 14792 2150
rect 14816 2148 14872 2150
rect 14896 2148 14952 2150
rect 14976 2148 15032 2150
<< metal3 >>
rect 1906 19072 2302 19073
rect 1906 19008 1912 19072
rect 1976 19008 1992 19072
rect 2056 19008 2072 19072
rect 2136 19008 2152 19072
rect 2216 19008 2232 19072
rect 2296 19008 2302 19072
rect 1906 19007 2302 19008
rect 7906 19072 8302 19073
rect 7906 19008 7912 19072
rect 7976 19008 7992 19072
rect 8056 19008 8072 19072
rect 8136 19008 8152 19072
rect 8216 19008 8232 19072
rect 8296 19008 8302 19072
rect 7906 19007 8302 19008
rect 13906 19072 14302 19073
rect 13906 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14152 19072
rect 14216 19008 14232 19072
rect 14296 19008 14302 19072
rect 13906 19007 14302 19008
rect 2646 18528 3042 18529
rect 2646 18464 2652 18528
rect 2716 18464 2732 18528
rect 2796 18464 2812 18528
rect 2876 18464 2892 18528
rect 2956 18464 2972 18528
rect 3036 18464 3042 18528
rect 2646 18463 3042 18464
rect 8646 18528 9042 18529
rect 8646 18464 8652 18528
rect 8716 18464 8732 18528
rect 8796 18464 8812 18528
rect 8876 18464 8892 18528
rect 8956 18464 8972 18528
rect 9036 18464 9042 18528
rect 8646 18463 9042 18464
rect 14646 18528 15042 18529
rect 14646 18464 14652 18528
rect 14716 18464 14732 18528
rect 14796 18464 14812 18528
rect 14876 18464 14892 18528
rect 14956 18464 14972 18528
rect 15036 18464 15042 18528
rect 14646 18463 15042 18464
rect 16665 18052 16731 18053
rect 16614 18050 16620 18052
rect 16574 17990 16620 18050
rect 16684 18048 16731 18052
rect 16726 17992 16731 18048
rect 16614 17988 16620 17990
rect 16684 17988 16731 17992
rect 16665 17987 16731 17988
rect 1906 17984 2302 17985
rect 1906 17920 1912 17984
rect 1976 17920 1992 17984
rect 2056 17920 2072 17984
rect 2136 17920 2152 17984
rect 2216 17920 2232 17984
rect 2296 17920 2302 17984
rect 1906 17919 2302 17920
rect 7906 17984 8302 17985
rect 7906 17920 7912 17984
rect 7976 17920 7992 17984
rect 8056 17920 8072 17984
rect 8136 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8302 17984
rect 7906 17919 8302 17920
rect 13906 17984 14302 17985
rect 13906 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14152 17984
rect 14216 17920 14232 17984
rect 14296 17920 14302 17984
rect 13906 17919 14302 17920
rect 2646 17440 3042 17441
rect 2646 17376 2652 17440
rect 2716 17376 2732 17440
rect 2796 17376 2812 17440
rect 2876 17376 2892 17440
rect 2956 17376 2972 17440
rect 3036 17376 3042 17440
rect 2646 17375 3042 17376
rect 8646 17440 9042 17441
rect 8646 17376 8652 17440
rect 8716 17376 8732 17440
rect 8796 17376 8812 17440
rect 8876 17376 8892 17440
rect 8956 17376 8972 17440
rect 9036 17376 9042 17440
rect 8646 17375 9042 17376
rect 14646 17440 15042 17441
rect 14646 17376 14652 17440
rect 14716 17376 14732 17440
rect 14796 17376 14812 17440
rect 14876 17376 14892 17440
rect 14956 17376 14972 17440
rect 15036 17376 15042 17440
rect 14646 17375 15042 17376
rect 1906 16896 2302 16897
rect 1906 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2302 16896
rect 1906 16831 2302 16832
rect 7906 16896 8302 16897
rect 7906 16832 7912 16896
rect 7976 16832 7992 16896
rect 8056 16832 8072 16896
rect 8136 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8302 16896
rect 7906 16831 8302 16832
rect 13906 16896 14302 16897
rect 13906 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14152 16896
rect 14216 16832 14232 16896
rect 14296 16832 14302 16896
rect 13906 16831 14302 16832
rect 2646 16352 3042 16353
rect 2646 16288 2652 16352
rect 2716 16288 2732 16352
rect 2796 16288 2812 16352
rect 2876 16288 2892 16352
rect 2956 16288 2972 16352
rect 3036 16288 3042 16352
rect 2646 16287 3042 16288
rect 8646 16352 9042 16353
rect 8646 16288 8652 16352
rect 8716 16288 8732 16352
rect 8796 16288 8812 16352
rect 8876 16288 8892 16352
rect 8956 16288 8972 16352
rect 9036 16288 9042 16352
rect 8646 16287 9042 16288
rect 14646 16352 15042 16353
rect 14646 16288 14652 16352
rect 14716 16288 14732 16352
rect 14796 16288 14812 16352
rect 14876 16288 14892 16352
rect 14956 16288 14972 16352
rect 15036 16288 15042 16352
rect 14646 16287 15042 16288
rect 0 15874 800 15904
rect 933 15874 999 15877
rect 0 15872 999 15874
rect 0 15816 938 15872
rect 994 15816 999 15872
rect 0 15814 999 15816
rect 0 15784 800 15814
rect 933 15811 999 15814
rect 1906 15808 2302 15809
rect 1906 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2302 15808
rect 1906 15743 2302 15744
rect 7906 15808 8302 15809
rect 7906 15744 7912 15808
rect 7976 15744 7992 15808
rect 8056 15744 8072 15808
rect 8136 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8302 15808
rect 7906 15743 8302 15744
rect 13906 15808 14302 15809
rect 13906 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14152 15808
rect 14216 15744 14232 15808
rect 14296 15744 14302 15808
rect 13906 15743 14302 15744
rect 2646 15264 3042 15265
rect 2646 15200 2652 15264
rect 2716 15200 2732 15264
rect 2796 15200 2812 15264
rect 2876 15200 2892 15264
rect 2956 15200 2972 15264
rect 3036 15200 3042 15264
rect 2646 15199 3042 15200
rect 8646 15264 9042 15265
rect 8646 15200 8652 15264
rect 8716 15200 8732 15264
rect 8796 15200 8812 15264
rect 8876 15200 8892 15264
rect 8956 15200 8972 15264
rect 9036 15200 9042 15264
rect 8646 15199 9042 15200
rect 14646 15264 15042 15265
rect 14646 15200 14652 15264
rect 14716 15200 14732 15264
rect 14796 15200 14812 15264
rect 14876 15200 14892 15264
rect 14956 15200 14972 15264
rect 15036 15200 15042 15264
rect 14646 15199 15042 15200
rect 1906 14720 2302 14721
rect 1906 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2302 14720
rect 1906 14655 2302 14656
rect 7906 14720 8302 14721
rect 7906 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8302 14720
rect 7906 14655 8302 14656
rect 13906 14720 14302 14721
rect 13906 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14302 14720
rect 13906 14655 14302 14656
rect 6361 14378 6427 14381
rect 8753 14378 8819 14381
rect 10041 14378 10107 14381
rect 13537 14378 13603 14381
rect 6361 14376 13603 14378
rect 6361 14320 6366 14376
rect 6422 14320 8758 14376
rect 8814 14320 10046 14376
rect 10102 14320 13542 14376
rect 13598 14320 13603 14376
rect 6361 14318 13603 14320
rect 6361 14315 6427 14318
rect 8753 14315 8819 14318
rect 10041 14315 10107 14318
rect 13537 14315 13603 14318
rect 2646 14176 3042 14177
rect 2646 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3042 14176
rect 2646 14111 3042 14112
rect 8646 14176 9042 14177
rect 8646 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9042 14176
rect 8646 14111 9042 14112
rect 14646 14176 15042 14177
rect 14646 14112 14652 14176
rect 14716 14112 14732 14176
rect 14796 14112 14812 14176
rect 14876 14112 14892 14176
rect 14956 14112 14972 14176
rect 15036 14112 15042 14176
rect 14646 14111 15042 14112
rect 1906 13632 2302 13633
rect 1906 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2302 13632
rect 1906 13567 2302 13568
rect 7906 13632 8302 13633
rect 7906 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8302 13632
rect 7906 13567 8302 13568
rect 13906 13632 14302 13633
rect 13906 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14302 13632
rect 13906 13567 14302 13568
rect 2646 13088 3042 13089
rect 2646 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3042 13088
rect 2646 13023 3042 13024
rect 8646 13088 9042 13089
rect 8646 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9042 13088
rect 8646 13023 9042 13024
rect 14646 13088 15042 13089
rect 14646 13024 14652 13088
rect 14716 13024 14732 13088
rect 14796 13024 14812 13088
rect 14876 13024 14892 13088
rect 14956 13024 14972 13088
rect 15036 13024 15042 13088
rect 14646 13023 15042 13024
rect 1906 12544 2302 12545
rect 1906 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2302 12544
rect 1906 12479 2302 12480
rect 7906 12544 8302 12545
rect 7906 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8302 12544
rect 7906 12479 8302 12480
rect 13906 12544 14302 12545
rect 13906 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14302 12544
rect 13906 12479 14302 12480
rect 2646 12000 3042 12001
rect 2646 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3042 12000
rect 2646 11935 3042 11936
rect 8646 12000 9042 12001
rect 8646 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9042 12000
rect 8646 11935 9042 11936
rect 14646 12000 15042 12001
rect 14646 11936 14652 12000
rect 14716 11936 14732 12000
rect 14796 11936 14812 12000
rect 14876 11936 14892 12000
rect 14956 11936 14972 12000
rect 15036 11936 15042 12000
rect 14646 11935 15042 11936
rect 1906 11456 2302 11457
rect 1906 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2302 11456
rect 1906 11391 2302 11392
rect 7906 11456 8302 11457
rect 7906 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8302 11456
rect 7906 11391 8302 11392
rect 13906 11456 14302 11457
rect 13906 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14302 11456
rect 13906 11391 14302 11392
rect 11329 11114 11395 11117
rect 11329 11112 16590 11114
rect 11329 11056 11334 11112
rect 11390 11056 16590 11112
rect 11329 11054 16590 11056
rect 11329 11051 11395 11054
rect 2646 10912 3042 10913
rect 2646 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3042 10912
rect 2646 10847 3042 10848
rect 8646 10912 9042 10913
rect 8646 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9042 10912
rect 8646 10847 9042 10848
rect 14646 10912 15042 10913
rect 14646 10848 14652 10912
rect 14716 10848 14732 10912
rect 14796 10848 14812 10912
rect 14876 10848 14892 10912
rect 14956 10848 14972 10912
rect 15036 10848 15042 10912
rect 14646 10847 15042 10848
rect 16530 10706 16590 11054
rect 18598 10706 19398 10736
rect 16530 10646 19398 10706
rect 18598 10616 19398 10646
rect 1906 10368 2302 10369
rect 1906 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2302 10368
rect 1906 10303 2302 10304
rect 7906 10368 8302 10369
rect 7906 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8302 10368
rect 7906 10303 8302 10304
rect 13906 10368 14302 10369
rect 13906 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14302 10368
rect 13906 10303 14302 10304
rect 2646 9824 3042 9825
rect 2646 9760 2652 9824
rect 2716 9760 2732 9824
rect 2796 9760 2812 9824
rect 2876 9760 2892 9824
rect 2956 9760 2972 9824
rect 3036 9760 3042 9824
rect 2646 9759 3042 9760
rect 8646 9824 9042 9825
rect 8646 9760 8652 9824
rect 8716 9760 8732 9824
rect 8796 9760 8812 9824
rect 8876 9760 8892 9824
rect 8956 9760 8972 9824
rect 9036 9760 9042 9824
rect 8646 9759 9042 9760
rect 14646 9824 15042 9825
rect 14646 9760 14652 9824
rect 14716 9760 14732 9824
rect 14796 9760 14812 9824
rect 14876 9760 14892 9824
rect 14956 9760 14972 9824
rect 15036 9760 15042 9824
rect 14646 9759 15042 9760
rect 1906 9280 2302 9281
rect 1906 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2302 9280
rect 1906 9215 2302 9216
rect 7906 9280 8302 9281
rect 7906 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8302 9280
rect 7906 9215 8302 9216
rect 13906 9280 14302 9281
rect 13906 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14152 9280
rect 14216 9216 14232 9280
rect 14296 9216 14302 9280
rect 13906 9215 14302 9216
rect 2646 8736 3042 8737
rect 2646 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3042 8736
rect 2646 8671 3042 8672
rect 8646 8736 9042 8737
rect 8646 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9042 8736
rect 8646 8671 9042 8672
rect 14646 8736 15042 8737
rect 14646 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15042 8736
rect 14646 8671 15042 8672
rect 5993 8530 6059 8533
rect 8753 8530 8819 8533
rect 9857 8530 9923 8533
rect 13813 8530 13879 8533
rect 14641 8530 14707 8533
rect 5993 8528 14707 8530
rect 5993 8472 5998 8528
rect 6054 8472 8758 8528
rect 8814 8472 9862 8528
rect 9918 8472 13818 8528
rect 13874 8472 14646 8528
rect 14702 8472 14707 8528
rect 5993 8470 14707 8472
rect 5993 8467 6059 8470
rect 8753 8467 8819 8470
rect 9857 8467 9923 8470
rect 13813 8467 13879 8470
rect 14641 8467 14707 8470
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 13906 8192 14302 8193
rect 13906 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14302 8192
rect 13906 8127 14302 8128
rect 2646 7648 3042 7649
rect 2646 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3042 7648
rect 2646 7583 3042 7584
rect 8646 7648 9042 7649
rect 8646 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9042 7648
rect 8646 7583 9042 7584
rect 14646 7648 15042 7649
rect 14646 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15042 7648
rect 14646 7583 15042 7584
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 13906 7104 14302 7105
rect 13906 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14302 7104
rect 13906 7039 14302 7040
rect 2646 6560 3042 6561
rect 2646 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3042 6560
rect 2646 6495 3042 6496
rect 8646 6560 9042 6561
rect 8646 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9042 6560
rect 8646 6495 9042 6496
rect 14646 6560 15042 6561
rect 14646 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15042 6560
rect 14646 6495 15042 6496
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 13906 6016 14302 6017
rect 13906 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14302 6016
rect 13906 5951 14302 5952
rect 16573 5812 16639 5813
rect 16573 5808 16620 5812
rect 16684 5810 16690 5812
rect 16573 5752 16578 5808
rect 16573 5748 16620 5752
rect 16684 5750 16730 5810
rect 16684 5748 16690 5750
rect 16573 5747 16639 5748
rect 2646 5472 3042 5473
rect 2646 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3042 5472
rect 2646 5407 3042 5408
rect 8646 5472 9042 5473
rect 8646 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9042 5472
rect 8646 5407 9042 5408
rect 14646 5472 15042 5473
rect 14646 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15042 5472
rect 14646 5407 15042 5408
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 13906 4928 14302 4929
rect 13906 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14302 4928
rect 13906 4863 14302 4864
rect 2646 4384 3042 4385
rect 2646 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3042 4384
rect 2646 4319 3042 4320
rect 8646 4384 9042 4385
rect 8646 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9042 4384
rect 8646 4319 9042 4320
rect 14646 4384 15042 4385
rect 14646 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15042 4384
rect 14646 4319 15042 4320
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 13906 3840 14302 3841
rect 13906 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14302 3840
rect 13906 3775 14302 3776
rect 2646 3296 3042 3297
rect 2646 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3042 3296
rect 2646 3231 3042 3232
rect 8646 3296 9042 3297
rect 8646 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9042 3296
rect 8646 3231 9042 3232
rect 14646 3296 15042 3297
rect 14646 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15042 3296
rect 14646 3231 15042 3232
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 13906 2752 14302 2753
rect 13906 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14302 2752
rect 13906 2687 14302 2688
rect 2646 2208 3042 2209
rect 2646 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3042 2208
rect 2646 2143 3042 2144
rect 8646 2208 9042 2209
rect 8646 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9042 2208
rect 8646 2143 9042 2144
rect 14646 2208 15042 2209
rect 14646 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15042 2208
rect 14646 2143 15042 2144
<< via3 >>
rect 1912 19068 1976 19072
rect 1912 19012 1916 19068
rect 1916 19012 1972 19068
rect 1972 19012 1976 19068
rect 1912 19008 1976 19012
rect 1992 19068 2056 19072
rect 1992 19012 1996 19068
rect 1996 19012 2052 19068
rect 2052 19012 2056 19068
rect 1992 19008 2056 19012
rect 2072 19068 2136 19072
rect 2072 19012 2076 19068
rect 2076 19012 2132 19068
rect 2132 19012 2136 19068
rect 2072 19008 2136 19012
rect 2152 19068 2216 19072
rect 2152 19012 2156 19068
rect 2156 19012 2212 19068
rect 2212 19012 2216 19068
rect 2152 19008 2216 19012
rect 2232 19068 2296 19072
rect 2232 19012 2236 19068
rect 2236 19012 2292 19068
rect 2292 19012 2296 19068
rect 2232 19008 2296 19012
rect 7912 19068 7976 19072
rect 7912 19012 7916 19068
rect 7916 19012 7972 19068
rect 7972 19012 7976 19068
rect 7912 19008 7976 19012
rect 7992 19068 8056 19072
rect 7992 19012 7996 19068
rect 7996 19012 8052 19068
rect 8052 19012 8056 19068
rect 7992 19008 8056 19012
rect 8072 19068 8136 19072
rect 8072 19012 8076 19068
rect 8076 19012 8132 19068
rect 8132 19012 8136 19068
rect 8072 19008 8136 19012
rect 8152 19068 8216 19072
rect 8152 19012 8156 19068
rect 8156 19012 8212 19068
rect 8212 19012 8216 19068
rect 8152 19008 8216 19012
rect 8232 19068 8296 19072
rect 8232 19012 8236 19068
rect 8236 19012 8292 19068
rect 8292 19012 8296 19068
rect 8232 19008 8296 19012
rect 13912 19068 13976 19072
rect 13912 19012 13916 19068
rect 13916 19012 13972 19068
rect 13972 19012 13976 19068
rect 13912 19008 13976 19012
rect 13992 19068 14056 19072
rect 13992 19012 13996 19068
rect 13996 19012 14052 19068
rect 14052 19012 14056 19068
rect 13992 19008 14056 19012
rect 14072 19068 14136 19072
rect 14072 19012 14076 19068
rect 14076 19012 14132 19068
rect 14132 19012 14136 19068
rect 14072 19008 14136 19012
rect 14152 19068 14216 19072
rect 14152 19012 14156 19068
rect 14156 19012 14212 19068
rect 14212 19012 14216 19068
rect 14152 19008 14216 19012
rect 14232 19068 14296 19072
rect 14232 19012 14236 19068
rect 14236 19012 14292 19068
rect 14292 19012 14296 19068
rect 14232 19008 14296 19012
rect 2652 18524 2716 18528
rect 2652 18468 2656 18524
rect 2656 18468 2712 18524
rect 2712 18468 2716 18524
rect 2652 18464 2716 18468
rect 2732 18524 2796 18528
rect 2732 18468 2736 18524
rect 2736 18468 2792 18524
rect 2792 18468 2796 18524
rect 2732 18464 2796 18468
rect 2812 18524 2876 18528
rect 2812 18468 2816 18524
rect 2816 18468 2872 18524
rect 2872 18468 2876 18524
rect 2812 18464 2876 18468
rect 2892 18524 2956 18528
rect 2892 18468 2896 18524
rect 2896 18468 2952 18524
rect 2952 18468 2956 18524
rect 2892 18464 2956 18468
rect 2972 18524 3036 18528
rect 2972 18468 2976 18524
rect 2976 18468 3032 18524
rect 3032 18468 3036 18524
rect 2972 18464 3036 18468
rect 8652 18524 8716 18528
rect 8652 18468 8656 18524
rect 8656 18468 8712 18524
rect 8712 18468 8716 18524
rect 8652 18464 8716 18468
rect 8732 18524 8796 18528
rect 8732 18468 8736 18524
rect 8736 18468 8792 18524
rect 8792 18468 8796 18524
rect 8732 18464 8796 18468
rect 8812 18524 8876 18528
rect 8812 18468 8816 18524
rect 8816 18468 8872 18524
rect 8872 18468 8876 18524
rect 8812 18464 8876 18468
rect 8892 18524 8956 18528
rect 8892 18468 8896 18524
rect 8896 18468 8952 18524
rect 8952 18468 8956 18524
rect 8892 18464 8956 18468
rect 8972 18524 9036 18528
rect 8972 18468 8976 18524
rect 8976 18468 9032 18524
rect 9032 18468 9036 18524
rect 8972 18464 9036 18468
rect 14652 18524 14716 18528
rect 14652 18468 14656 18524
rect 14656 18468 14712 18524
rect 14712 18468 14716 18524
rect 14652 18464 14716 18468
rect 14732 18524 14796 18528
rect 14732 18468 14736 18524
rect 14736 18468 14792 18524
rect 14792 18468 14796 18524
rect 14732 18464 14796 18468
rect 14812 18524 14876 18528
rect 14812 18468 14816 18524
rect 14816 18468 14872 18524
rect 14872 18468 14876 18524
rect 14812 18464 14876 18468
rect 14892 18524 14956 18528
rect 14892 18468 14896 18524
rect 14896 18468 14952 18524
rect 14952 18468 14956 18524
rect 14892 18464 14956 18468
rect 14972 18524 15036 18528
rect 14972 18468 14976 18524
rect 14976 18468 15032 18524
rect 15032 18468 15036 18524
rect 14972 18464 15036 18468
rect 16620 18048 16684 18052
rect 16620 17992 16670 18048
rect 16670 17992 16684 18048
rect 16620 17988 16684 17992
rect 1912 17980 1976 17984
rect 1912 17924 1916 17980
rect 1916 17924 1972 17980
rect 1972 17924 1976 17980
rect 1912 17920 1976 17924
rect 1992 17980 2056 17984
rect 1992 17924 1996 17980
rect 1996 17924 2052 17980
rect 2052 17924 2056 17980
rect 1992 17920 2056 17924
rect 2072 17980 2136 17984
rect 2072 17924 2076 17980
rect 2076 17924 2132 17980
rect 2132 17924 2136 17980
rect 2072 17920 2136 17924
rect 2152 17980 2216 17984
rect 2152 17924 2156 17980
rect 2156 17924 2212 17980
rect 2212 17924 2216 17980
rect 2152 17920 2216 17924
rect 2232 17980 2296 17984
rect 2232 17924 2236 17980
rect 2236 17924 2292 17980
rect 2292 17924 2296 17980
rect 2232 17920 2296 17924
rect 7912 17980 7976 17984
rect 7912 17924 7916 17980
rect 7916 17924 7972 17980
rect 7972 17924 7976 17980
rect 7912 17920 7976 17924
rect 7992 17980 8056 17984
rect 7992 17924 7996 17980
rect 7996 17924 8052 17980
rect 8052 17924 8056 17980
rect 7992 17920 8056 17924
rect 8072 17980 8136 17984
rect 8072 17924 8076 17980
rect 8076 17924 8132 17980
rect 8132 17924 8136 17980
rect 8072 17920 8136 17924
rect 8152 17980 8216 17984
rect 8152 17924 8156 17980
rect 8156 17924 8212 17980
rect 8212 17924 8216 17980
rect 8152 17920 8216 17924
rect 8232 17980 8296 17984
rect 8232 17924 8236 17980
rect 8236 17924 8292 17980
rect 8292 17924 8296 17980
rect 8232 17920 8296 17924
rect 13912 17980 13976 17984
rect 13912 17924 13916 17980
rect 13916 17924 13972 17980
rect 13972 17924 13976 17980
rect 13912 17920 13976 17924
rect 13992 17980 14056 17984
rect 13992 17924 13996 17980
rect 13996 17924 14052 17980
rect 14052 17924 14056 17980
rect 13992 17920 14056 17924
rect 14072 17980 14136 17984
rect 14072 17924 14076 17980
rect 14076 17924 14132 17980
rect 14132 17924 14136 17980
rect 14072 17920 14136 17924
rect 14152 17980 14216 17984
rect 14152 17924 14156 17980
rect 14156 17924 14212 17980
rect 14212 17924 14216 17980
rect 14152 17920 14216 17924
rect 14232 17980 14296 17984
rect 14232 17924 14236 17980
rect 14236 17924 14292 17980
rect 14292 17924 14296 17980
rect 14232 17920 14296 17924
rect 2652 17436 2716 17440
rect 2652 17380 2656 17436
rect 2656 17380 2712 17436
rect 2712 17380 2716 17436
rect 2652 17376 2716 17380
rect 2732 17436 2796 17440
rect 2732 17380 2736 17436
rect 2736 17380 2792 17436
rect 2792 17380 2796 17436
rect 2732 17376 2796 17380
rect 2812 17436 2876 17440
rect 2812 17380 2816 17436
rect 2816 17380 2872 17436
rect 2872 17380 2876 17436
rect 2812 17376 2876 17380
rect 2892 17436 2956 17440
rect 2892 17380 2896 17436
rect 2896 17380 2952 17436
rect 2952 17380 2956 17436
rect 2892 17376 2956 17380
rect 2972 17436 3036 17440
rect 2972 17380 2976 17436
rect 2976 17380 3032 17436
rect 3032 17380 3036 17436
rect 2972 17376 3036 17380
rect 8652 17436 8716 17440
rect 8652 17380 8656 17436
rect 8656 17380 8712 17436
rect 8712 17380 8716 17436
rect 8652 17376 8716 17380
rect 8732 17436 8796 17440
rect 8732 17380 8736 17436
rect 8736 17380 8792 17436
rect 8792 17380 8796 17436
rect 8732 17376 8796 17380
rect 8812 17436 8876 17440
rect 8812 17380 8816 17436
rect 8816 17380 8872 17436
rect 8872 17380 8876 17436
rect 8812 17376 8876 17380
rect 8892 17436 8956 17440
rect 8892 17380 8896 17436
rect 8896 17380 8952 17436
rect 8952 17380 8956 17436
rect 8892 17376 8956 17380
rect 8972 17436 9036 17440
rect 8972 17380 8976 17436
rect 8976 17380 9032 17436
rect 9032 17380 9036 17436
rect 8972 17376 9036 17380
rect 14652 17436 14716 17440
rect 14652 17380 14656 17436
rect 14656 17380 14712 17436
rect 14712 17380 14716 17436
rect 14652 17376 14716 17380
rect 14732 17436 14796 17440
rect 14732 17380 14736 17436
rect 14736 17380 14792 17436
rect 14792 17380 14796 17436
rect 14732 17376 14796 17380
rect 14812 17436 14876 17440
rect 14812 17380 14816 17436
rect 14816 17380 14872 17436
rect 14872 17380 14876 17436
rect 14812 17376 14876 17380
rect 14892 17436 14956 17440
rect 14892 17380 14896 17436
rect 14896 17380 14952 17436
rect 14952 17380 14956 17436
rect 14892 17376 14956 17380
rect 14972 17436 15036 17440
rect 14972 17380 14976 17436
rect 14976 17380 15032 17436
rect 15032 17380 15036 17436
rect 14972 17376 15036 17380
rect 1912 16892 1976 16896
rect 1912 16836 1916 16892
rect 1916 16836 1972 16892
rect 1972 16836 1976 16892
rect 1912 16832 1976 16836
rect 1992 16892 2056 16896
rect 1992 16836 1996 16892
rect 1996 16836 2052 16892
rect 2052 16836 2056 16892
rect 1992 16832 2056 16836
rect 2072 16892 2136 16896
rect 2072 16836 2076 16892
rect 2076 16836 2132 16892
rect 2132 16836 2136 16892
rect 2072 16832 2136 16836
rect 2152 16892 2216 16896
rect 2152 16836 2156 16892
rect 2156 16836 2212 16892
rect 2212 16836 2216 16892
rect 2152 16832 2216 16836
rect 2232 16892 2296 16896
rect 2232 16836 2236 16892
rect 2236 16836 2292 16892
rect 2292 16836 2296 16892
rect 2232 16832 2296 16836
rect 7912 16892 7976 16896
rect 7912 16836 7916 16892
rect 7916 16836 7972 16892
rect 7972 16836 7976 16892
rect 7912 16832 7976 16836
rect 7992 16892 8056 16896
rect 7992 16836 7996 16892
rect 7996 16836 8052 16892
rect 8052 16836 8056 16892
rect 7992 16832 8056 16836
rect 8072 16892 8136 16896
rect 8072 16836 8076 16892
rect 8076 16836 8132 16892
rect 8132 16836 8136 16892
rect 8072 16832 8136 16836
rect 8152 16892 8216 16896
rect 8152 16836 8156 16892
rect 8156 16836 8212 16892
rect 8212 16836 8216 16892
rect 8152 16832 8216 16836
rect 8232 16892 8296 16896
rect 8232 16836 8236 16892
rect 8236 16836 8292 16892
rect 8292 16836 8296 16892
rect 8232 16832 8296 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 14152 16892 14216 16896
rect 14152 16836 14156 16892
rect 14156 16836 14212 16892
rect 14212 16836 14216 16892
rect 14152 16832 14216 16836
rect 14232 16892 14296 16896
rect 14232 16836 14236 16892
rect 14236 16836 14292 16892
rect 14292 16836 14296 16892
rect 14232 16832 14296 16836
rect 2652 16348 2716 16352
rect 2652 16292 2656 16348
rect 2656 16292 2712 16348
rect 2712 16292 2716 16348
rect 2652 16288 2716 16292
rect 2732 16348 2796 16352
rect 2732 16292 2736 16348
rect 2736 16292 2792 16348
rect 2792 16292 2796 16348
rect 2732 16288 2796 16292
rect 2812 16348 2876 16352
rect 2812 16292 2816 16348
rect 2816 16292 2872 16348
rect 2872 16292 2876 16348
rect 2812 16288 2876 16292
rect 2892 16348 2956 16352
rect 2892 16292 2896 16348
rect 2896 16292 2952 16348
rect 2952 16292 2956 16348
rect 2892 16288 2956 16292
rect 2972 16348 3036 16352
rect 2972 16292 2976 16348
rect 2976 16292 3032 16348
rect 3032 16292 3036 16348
rect 2972 16288 3036 16292
rect 8652 16348 8716 16352
rect 8652 16292 8656 16348
rect 8656 16292 8712 16348
rect 8712 16292 8716 16348
rect 8652 16288 8716 16292
rect 8732 16348 8796 16352
rect 8732 16292 8736 16348
rect 8736 16292 8792 16348
rect 8792 16292 8796 16348
rect 8732 16288 8796 16292
rect 8812 16348 8876 16352
rect 8812 16292 8816 16348
rect 8816 16292 8872 16348
rect 8872 16292 8876 16348
rect 8812 16288 8876 16292
rect 8892 16348 8956 16352
rect 8892 16292 8896 16348
rect 8896 16292 8952 16348
rect 8952 16292 8956 16348
rect 8892 16288 8956 16292
rect 8972 16348 9036 16352
rect 8972 16292 8976 16348
rect 8976 16292 9032 16348
rect 9032 16292 9036 16348
rect 8972 16288 9036 16292
rect 14652 16348 14716 16352
rect 14652 16292 14656 16348
rect 14656 16292 14712 16348
rect 14712 16292 14716 16348
rect 14652 16288 14716 16292
rect 14732 16348 14796 16352
rect 14732 16292 14736 16348
rect 14736 16292 14792 16348
rect 14792 16292 14796 16348
rect 14732 16288 14796 16292
rect 14812 16348 14876 16352
rect 14812 16292 14816 16348
rect 14816 16292 14872 16348
rect 14872 16292 14876 16348
rect 14812 16288 14876 16292
rect 14892 16348 14956 16352
rect 14892 16292 14896 16348
rect 14896 16292 14952 16348
rect 14952 16292 14956 16348
rect 14892 16288 14956 16292
rect 14972 16348 15036 16352
rect 14972 16292 14976 16348
rect 14976 16292 15032 16348
rect 15032 16292 15036 16348
rect 14972 16288 15036 16292
rect 1912 15804 1976 15808
rect 1912 15748 1916 15804
rect 1916 15748 1972 15804
rect 1972 15748 1976 15804
rect 1912 15744 1976 15748
rect 1992 15804 2056 15808
rect 1992 15748 1996 15804
rect 1996 15748 2052 15804
rect 2052 15748 2056 15804
rect 1992 15744 2056 15748
rect 2072 15804 2136 15808
rect 2072 15748 2076 15804
rect 2076 15748 2132 15804
rect 2132 15748 2136 15804
rect 2072 15744 2136 15748
rect 2152 15804 2216 15808
rect 2152 15748 2156 15804
rect 2156 15748 2212 15804
rect 2212 15748 2216 15804
rect 2152 15744 2216 15748
rect 2232 15804 2296 15808
rect 2232 15748 2236 15804
rect 2236 15748 2292 15804
rect 2292 15748 2296 15804
rect 2232 15744 2296 15748
rect 7912 15804 7976 15808
rect 7912 15748 7916 15804
rect 7916 15748 7972 15804
rect 7972 15748 7976 15804
rect 7912 15744 7976 15748
rect 7992 15804 8056 15808
rect 7992 15748 7996 15804
rect 7996 15748 8052 15804
rect 8052 15748 8056 15804
rect 7992 15744 8056 15748
rect 8072 15804 8136 15808
rect 8072 15748 8076 15804
rect 8076 15748 8132 15804
rect 8132 15748 8136 15804
rect 8072 15744 8136 15748
rect 8152 15804 8216 15808
rect 8152 15748 8156 15804
rect 8156 15748 8212 15804
rect 8212 15748 8216 15804
rect 8152 15744 8216 15748
rect 8232 15804 8296 15808
rect 8232 15748 8236 15804
rect 8236 15748 8292 15804
rect 8292 15748 8296 15804
rect 8232 15744 8296 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 14152 15804 14216 15808
rect 14152 15748 14156 15804
rect 14156 15748 14212 15804
rect 14212 15748 14216 15804
rect 14152 15744 14216 15748
rect 14232 15804 14296 15808
rect 14232 15748 14236 15804
rect 14236 15748 14292 15804
rect 14292 15748 14296 15804
rect 14232 15744 14296 15748
rect 2652 15260 2716 15264
rect 2652 15204 2656 15260
rect 2656 15204 2712 15260
rect 2712 15204 2716 15260
rect 2652 15200 2716 15204
rect 2732 15260 2796 15264
rect 2732 15204 2736 15260
rect 2736 15204 2792 15260
rect 2792 15204 2796 15260
rect 2732 15200 2796 15204
rect 2812 15260 2876 15264
rect 2812 15204 2816 15260
rect 2816 15204 2872 15260
rect 2872 15204 2876 15260
rect 2812 15200 2876 15204
rect 2892 15260 2956 15264
rect 2892 15204 2896 15260
rect 2896 15204 2952 15260
rect 2952 15204 2956 15260
rect 2892 15200 2956 15204
rect 2972 15260 3036 15264
rect 2972 15204 2976 15260
rect 2976 15204 3032 15260
rect 3032 15204 3036 15260
rect 2972 15200 3036 15204
rect 8652 15260 8716 15264
rect 8652 15204 8656 15260
rect 8656 15204 8712 15260
rect 8712 15204 8716 15260
rect 8652 15200 8716 15204
rect 8732 15260 8796 15264
rect 8732 15204 8736 15260
rect 8736 15204 8792 15260
rect 8792 15204 8796 15260
rect 8732 15200 8796 15204
rect 8812 15260 8876 15264
rect 8812 15204 8816 15260
rect 8816 15204 8872 15260
rect 8872 15204 8876 15260
rect 8812 15200 8876 15204
rect 8892 15260 8956 15264
rect 8892 15204 8896 15260
rect 8896 15204 8952 15260
rect 8952 15204 8956 15260
rect 8892 15200 8956 15204
rect 8972 15260 9036 15264
rect 8972 15204 8976 15260
rect 8976 15204 9032 15260
rect 9032 15204 9036 15260
rect 8972 15200 9036 15204
rect 14652 15260 14716 15264
rect 14652 15204 14656 15260
rect 14656 15204 14712 15260
rect 14712 15204 14716 15260
rect 14652 15200 14716 15204
rect 14732 15260 14796 15264
rect 14732 15204 14736 15260
rect 14736 15204 14792 15260
rect 14792 15204 14796 15260
rect 14732 15200 14796 15204
rect 14812 15260 14876 15264
rect 14812 15204 14816 15260
rect 14816 15204 14872 15260
rect 14872 15204 14876 15260
rect 14812 15200 14876 15204
rect 14892 15260 14956 15264
rect 14892 15204 14896 15260
rect 14896 15204 14952 15260
rect 14952 15204 14956 15260
rect 14892 15200 14956 15204
rect 14972 15260 15036 15264
rect 14972 15204 14976 15260
rect 14976 15204 15032 15260
rect 15032 15204 15036 15260
rect 14972 15200 15036 15204
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 7912 14716 7976 14720
rect 7912 14660 7916 14716
rect 7916 14660 7972 14716
rect 7972 14660 7976 14716
rect 7912 14656 7976 14660
rect 7992 14716 8056 14720
rect 7992 14660 7996 14716
rect 7996 14660 8052 14716
rect 8052 14660 8056 14716
rect 7992 14656 8056 14660
rect 8072 14716 8136 14720
rect 8072 14660 8076 14716
rect 8076 14660 8132 14716
rect 8132 14660 8136 14716
rect 8072 14656 8136 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 14152 14716 14216 14720
rect 14152 14660 14156 14716
rect 14156 14660 14212 14716
rect 14212 14660 14216 14716
rect 14152 14656 14216 14660
rect 14232 14716 14296 14720
rect 14232 14660 14236 14716
rect 14236 14660 14292 14716
rect 14292 14660 14296 14716
rect 14232 14656 14296 14660
rect 2652 14172 2716 14176
rect 2652 14116 2656 14172
rect 2656 14116 2712 14172
rect 2712 14116 2716 14172
rect 2652 14112 2716 14116
rect 2732 14172 2796 14176
rect 2732 14116 2736 14172
rect 2736 14116 2792 14172
rect 2792 14116 2796 14172
rect 2732 14112 2796 14116
rect 2812 14172 2876 14176
rect 2812 14116 2816 14172
rect 2816 14116 2872 14172
rect 2872 14116 2876 14172
rect 2812 14112 2876 14116
rect 2892 14172 2956 14176
rect 2892 14116 2896 14172
rect 2896 14116 2952 14172
rect 2952 14116 2956 14172
rect 2892 14112 2956 14116
rect 2972 14172 3036 14176
rect 2972 14116 2976 14172
rect 2976 14116 3032 14172
rect 3032 14116 3036 14172
rect 2972 14112 3036 14116
rect 8652 14172 8716 14176
rect 8652 14116 8656 14172
rect 8656 14116 8712 14172
rect 8712 14116 8716 14172
rect 8652 14112 8716 14116
rect 8732 14172 8796 14176
rect 8732 14116 8736 14172
rect 8736 14116 8792 14172
rect 8792 14116 8796 14172
rect 8732 14112 8796 14116
rect 8812 14172 8876 14176
rect 8812 14116 8816 14172
rect 8816 14116 8872 14172
rect 8872 14116 8876 14172
rect 8812 14112 8876 14116
rect 8892 14172 8956 14176
rect 8892 14116 8896 14172
rect 8896 14116 8952 14172
rect 8952 14116 8956 14172
rect 8892 14112 8956 14116
rect 8972 14172 9036 14176
rect 8972 14116 8976 14172
rect 8976 14116 9032 14172
rect 9032 14116 9036 14172
rect 8972 14112 9036 14116
rect 14652 14172 14716 14176
rect 14652 14116 14656 14172
rect 14656 14116 14712 14172
rect 14712 14116 14716 14172
rect 14652 14112 14716 14116
rect 14732 14172 14796 14176
rect 14732 14116 14736 14172
rect 14736 14116 14792 14172
rect 14792 14116 14796 14172
rect 14732 14112 14796 14116
rect 14812 14172 14876 14176
rect 14812 14116 14816 14172
rect 14816 14116 14872 14172
rect 14872 14116 14876 14172
rect 14812 14112 14876 14116
rect 14892 14172 14956 14176
rect 14892 14116 14896 14172
rect 14896 14116 14952 14172
rect 14952 14116 14956 14172
rect 14892 14112 14956 14116
rect 14972 14172 15036 14176
rect 14972 14116 14976 14172
rect 14976 14116 15032 14172
rect 15032 14116 15036 14172
rect 14972 14112 15036 14116
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 7912 13628 7976 13632
rect 7912 13572 7916 13628
rect 7916 13572 7972 13628
rect 7972 13572 7976 13628
rect 7912 13568 7976 13572
rect 7992 13628 8056 13632
rect 7992 13572 7996 13628
rect 7996 13572 8052 13628
rect 8052 13572 8056 13628
rect 7992 13568 8056 13572
rect 8072 13628 8136 13632
rect 8072 13572 8076 13628
rect 8076 13572 8132 13628
rect 8132 13572 8136 13628
rect 8072 13568 8136 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 14152 13628 14216 13632
rect 14152 13572 14156 13628
rect 14156 13572 14212 13628
rect 14212 13572 14216 13628
rect 14152 13568 14216 13572
rect 14232 13628 14296 13632
rect 14232 13572 14236 13628
rect 14236 13572 14292 13628
rect 14292 13572 14296 13628
rect 14232 13568 14296 13572
rect 2652 13084 2716 13088
rect 2652 13028 2656 13084
rect 2656 13028 2712 13084
rect 2712 13028 2716 13084
rect 2652 13024 2716 13028
rect 2732 13084 2796 13088
rect 2732 13028 2736 13084
rect 2736 13028 2792 13084
rect 2792 13028 2796 13084
rect 2732 13024 2796 13028
rect 2812 13084 2876 13088
rect 2812 13028 2816 13084
rect 2816 13028 2872 13084
rect 2872 13028 2876 13084
rect 2812 13024 2876 13028
rect 2892 13084 2956 13088
rect 2892 13028 2896 13084
rect 2896 13028 2952 13084
rect 2952 13028 2956 13084
rect 2892 13024 2956 13028
rect 2972 13084 3036 13088
rect 2972 13028 2976 13084
rect 2976 13028 3032 13084
rect 3032 13028 3036 13084
rect 2972 13024 3036 13028
rect 8652 13084 8716 13088
rect 8652 13028 8656 13084
rect 8656 13028 8712 13084
rect 8712 13028 8716 13084
rect 8652 13024 8716 13028
rect 8732 13084 8796 13088
rect 8732 13028 8736 13084
rect 8736 13028 8792 13084
rect 8792 13028 8796 13084
rect 8732 13024 8796 13028
rect 8812 13084 8876 13088
rect 8812 13028 8816 13084
rect 8816 13028 8872 13084
rect 8872 13028 8876 13084
rect 8812 13024 8876 13028
rect 8892 13084 8956 13088
rect 8892 13028 8896 13084
rect 8896 13028 8952 13084
rect 8952 13028 8956 13084
rect 8892 13024 8956 13028
rect 8972 13084 9036 13088
rect 8972 13028 8976 13084
rect 8976 13028 9032 13084
rect 9032 13028 9036 13084
rect 8972 13024 9036 13028
rect 14652 13084 14716 13088
rect 14652 13028 14656 13084
rect 14656 13028 14712 13084
rect 14712 13028 14716 13084
rect 14652 13024 14716 13028
rect 14732 13084 14796 13088
rect 14732 13028 14736 13084
rect 14736 13028 14792 13084
rect 14792 13028 14796 13084
rect 14732 13024 14796 13028
rect 14812 13084 14876 13088
rect 14812 13028 14816 13084
rect 14816 13028 14872 13084
rect 14872 13028 14876 13084
rect 14812 13024 14876 13028
rect 14892 13084 14956 13088
rect 14892 13028 14896 13084
rect 14896 13028 14952 13084
rect 14952 13028 14956 13084
rect 14892 13024 14956 13028
rect 14972 13084 15036 13088
rect 14972 13028 14976 13084
rect 14976 13028 15032 13084
rect 15032 13028 15036 13084
rect 14972 13024 15036 13028
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 7912 12540 7976 12544
rect 7912 12484 7916 12540
rect 7916 12484 7972 12540
rect 7972 12484 7976 12540
rect 7912 12480 7976 12484
rect 7992 12540 8056 12544
rect 7992 12484 7996 12540
rect 7996 12484 8052 12540
rect 8052 12484 8056 12540
rect 7992 12480 8056 12484
rect 8072 12540 8136 12544
rect 8072 12484 8076 12540
rect 8076 12484 8132 12540
rect 8132 12484 8136 12540
rect 8072 12480 8136 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 14152 12540 14216 12544
rect 14152 12484 14156 12540
rect 14156 12484 14212 12540
rect 14212 12484 14216 12540
rect 14152 12480 14216 12484
rect 14232 12540 14296 12544
rect 14232 12484 14236 12540
rect 14236 12484 14292 12540
rect 14292 12484 14296 12540
rect 14232 12480 14296 12484
rect 2652 11996 2716 12000
rect 2652 11940 2656 11996
rect 2656 11940 2712 11996
rect 2712 11940 2716 11996
rect 2652 11936 2716 11940
rect 2732 11996 2796 12000
rect 2732 11940 2736 11996
rect 2736 11940 2792 11996
rect 2792 11940 2796 11996
rect 2732 11936 2796 11940
rect 2812 11996 2876 12000
rect 2812 11940 2816 11996
rect 2816 11940 2872 11996
rect 2872 11940 2876 11996
rect 2812 11936 2876 11940
rect 2892 11996 2956 12000
rect 2892 11940 2896 11996
rect 2896 11940 2952 11996
rect 2952 11940 2956 11996
rect 2892 11936 2956 11940
rect 2972 11996 3036 12000
rect 2972 11940 2976 11996
rect 2976 11940 3032 11996
rect 3032 11940 3036 11996
rect 2972 11936 3036 11940
rect 8652 11996 8716 12000
rect 8652 11940 8656 11996
rect 8656 11940 8712 11996
rect 8712 11940 8716 11996
rect 8652 11936 8716 11940
rect 8732 11996 8796 12000
rect 8732 11940 8736 11996
rect 8736 11940 8792 11996
rect 8792 11940 8796 11996
rect 8732 11936 8796 11940
rect 8812 11996 8876 12000
rect 8812 11940 8816 11996
rect 8816 11940 8872 11996
rect 8872 11940 8876 11996
rect 8812 11936 8876 11940
rect 8892 11996 8956 12000
rect 8892 11940 8896 11996
rect 8896 11940 8952 11996
rect 8952 11940 8956 11996
rect 8892 11936 8956 11940
rect 8972 11996 9036 12000
rect 8972 11940 8976 11996
rect 8976 11940 9032 11996
rect 9032 11940 9036 11996
rect 8972 11936 9036 11940
rect 14652 11996 14716 12000
rect 14652 11940 14656 11996
rect 14656 11940 14712 11996
rect 14712 11940 14716 11996
rect 14652 11936 14716 11940
rect 14732 11996 14796 12000
rect 14732 11940 14736 11996
rect 14736 11940 14792 11996
rect 14792 11940 14796 11996
rect 14732 11936 14796 11940
rect 14812 11996 14876 12000
rect 14812 11940 14816 11996
rect 14816 11940 14872 11996
rect 14872 11940 14876 11996
rect 14812 11936 14876 11940
rect 14892 11996 14956 12000
rect 14892 11940 14896 11996
rect 14896 11940 14952 11996
rect 14952 11940 14956 11996
rect 14892 11936 14956 11940
rect 14972 11996 15036 12000
rect 14972 11940 14976 11996
rect 14976 11940 15032 11996
rect 15032 11940 15036 11996
rect 14972 11936 15036 11940
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 7912 11452 7976 11456
rect 7912 11396 7916 11452
rect 7916 11396 7972 11452
rect 7972 11396 7976 11452
rect 7912 11392 7976 11396
rect 7992 11452 8056 11456
rect 7992 11396 7996 11452
rect 7996 11396 8052 11452
rect 8052 11396 8056 11452
rect 7992 11392 8056 11396
rect 8072 11452 8136 11456
rect 8072 11396 8076 11452
rect 8076 11396 8132 11452
rect 8132 11396 8136 11452
rect 8072 11392 8136 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 14152 11452 14216 11456
rect 14152 11396 14156 11452
rect 14156 11396 14212 11452
rect 14212 11396 14216 11452
rect 14152 11392 14216 11396
rect 14232 11452 14296 11456
rect 14232 11396 14236 11452
rect 14236 11396 14292 11452
rect 14292 11396 14296 11452
rect 14232 11392 14296 11396
rect 2652 10908 2716 10912
rect 2652 10852 2656 10908
rect 2656 10852 2712 10908
rect 2712 10852 2716 10908
rect 2652 10848 2716 10852
rect 2732 10908 2796 10912
rect 2732 10852 2736 10908
rect 2736 10852 2792 10908
rect 2792 10852 2796 10908
rect 2732 10848 2796 10852
rect 2812 10908 2876 10912
rect 2812 10852 2816 10908
rect 2816 10852 2872 10908
rect 2872 10852 2876 10908
rect 2812 10848 2876 10852
rect 2892 10908 2956 10912
rect 2892 10852 2896 10908
rect 2896 10852 2952 10908
rect 2952 10852 2956 10908
rect 2892 10848 2956 10852
rect 2972 10908 3036 10912
rect 2972 10852 2976 10908
rect 2976 10852 3032 10908
rect 3032 10852 3036 10908
rect 2972 10848 3036 10852
rect 8652 10908 8716 10912
rect 8652 10852 8656 10908
rect 8656 10852 8712 10908
rect 8712 10852 8716 10908
rect 8652 10848 8716 10852
rect 8732 10908 8796 10912
rect 8732 10852 8736 10908
rect 8736 10852 8792 10908
rect 8792 10852 8796 10908
rect 8732 10848 8796 10852
rect 8812 10908 8876 10912
rect 8812 10852 8816 10908
rect 8816 10852 8872 10908
rect 8872 10852 8876 10908
rect 8812 10848 8876 10852
rect 8892 10908 8956 10912
rect 8892 10852 8896 10908
rect 8896 10852 8952 10908
rect 8952 10852 8956 10908
rect 8892 10848 8956 10852
rect 8972 10908 9036 10912
rect 8972 10852 8976 10908
rect 8976 10852 9032 10908
rect 9032 10852 9036 10908
rect 8972 10848 9036 10852
rect 14652 10908 14716 10912
rect 14652 10852 14656 10908
rect 14656 10852 14712 10908
rect 14712 10852 14716 10908
rect 14652 10848 14716 10852
rect 14732 10908 14796 10912
rect 14732 10852 14736 10908
rect 14736 10852 14792 10908
rect 14792 10852 14796 10908
rect 14732 10848 14796 10852
rect 14812 10908 14876 10912
rect 14812 10852 14816 10908
rect 14816 10852 14872 10908
rect 14872 10852 14876 10908
rect 14812 10848 14876 10852
rect 14892 10908 14956 10912
rect 14892 10852 14896 10908
rect 14896 10852 14952 10908
rect 14952 10852 14956 10908
rect 14892 10848 14956 10852
rect 14972 10908 15036 10912
rect 14972 10852 14976 10908
rect 14976 10852 15032 10908
rect 15032 10852 15036 10908
rect 14972 10848 15036 10852
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 7912 10364 7976 10368
rect 7912 10308 7916 10364
rect 7916 10308 7972 10364
rect 7972 10308 7976 10364
rect 7912 10304 7976 10308
rect 7992 10364 8056 10368
rect 7992 10308 7996 10364
rect 7996 10308 8052 10364
rect 8052 10308 8056 10364
rect 7992 10304 8056 10308
rect 8072 10364 8136 10368
rect 8072 10308 8076 10364
rect 8076 10308 8132 10364
rect 8132 10308 8136 10364
rect 8072 10304 8136 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 14152 10364 14216 10368
rect 14152 10308 14156 10364
rect 14156 10308 14212 10364
rect 14212 10308 14216 10364
rect 14152 10304 14216 10308
rect 14232 10364 14296 10368
rect 14232 10308 14236 10364
rect 14236 10308 14292 10364
rect 14292 10308 14296 10364
rect 14232 10304 14296 10308
rect 2652 9820 2716 9824
rect 2652 9764 2656 9820
rect 2656 9764 2712 9820
rect 2712 9764 2716 9820
rect 2652 9760 2716 9764
rect 2732 9820 2796 9824
rect 2732 9764 2736 9820
rect 2736 9764 2792 9820
rect 2792 9764 2796 9820
rect 2732 9760 2796 9764
rect 2812 9820 2876 9824
rect 2812 9764 2816 9820
rect 2816 9764 2872 9820
rect 2872 9764 2876 9820
rect 2812 9760 2876 9764
rect 2892 9820 2956 9824
rect 2892 9764 2896 9820
rect 2896 9764 2952 9820
rect 2952 9764 2956 9820
rect 2892 9760 2956 9764
rect 2972 9820 3036 9824
rect 2972 9764 2976 9820
rect 2976 9764 3032 9820
rect 3032 9764 3036 9820
rect 2972 9760 3036 9764
rect 8652 9820 8716 9824
rect 8652 9764 8656 9820
rect 8656 9764 8712 9820
rect 8712 9764 8716 9820
rect 8652 9760 8716 9764
rect 8732 9820 8796 9824
rect 8732 9764 8736 9820
rect 8736 9764 8792 9820
rect 8792 9764 8796 9820
rect 8732 9760 8796 9764
rect 8812 9820 8876 9824
rect 8812 9764 8816 9820
rect 8816 9764 8872 9820
rect 8872 9764 8876 9820
rect 8812 9760 8876 9764
rect 8892 9820 8956 9824
rect 8892 9764 8896 9820
rect 8896 9764 8952 9820
rect 8952 9764 8956 9820
rect 8892 9760 8956 9764
rect 8972 9820 9036 9824
rect 8972 9764 8976 9820
rect 8976 9764 9032 9820
rect 9032 9764 9036 9820
rect 8972 9760 9036 9764
rect 14652 9820 14716 9824
rect 14652 9764 14656 9820
rect 14656 9764 14712 9820
rect 14712 9764 14716 9820
rect 14652 9760 14716 9764
rect 14732 9820 14796 9824
rect 14732 9764 14736 9820
rect 14736 9764 14792 9820
rect 14792 9764 14796 9820
rect 14732 9760 14796 9764
rect 14812 9820 14876 9824
rect 14812 9764 14816 9820
rect 14816 9764 14872 9820
rect 14872 9764 14876 9820
rect 14812 9760 14876 9764
rect 14892 9820 14956 9824
rect 14892 9764 14896 9820
rect 14896 9764 14952 9820
rect 14952 9764 14956 9820
rect 14892 9760 14956 9764
rect 14972 9820 15036 9824
rect 14972 9764 14976 9820
rect 14976 9764 15032 9820
rect 15032 9764 15036 9820
rect 14972 9760 15036 9764
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 8072 9276 8136 9280
rect 8072 9220 8076 9276
rect 8076 9220 8132 9276
rect 8132 9220 8136 9276
rect 8072 9216 8136 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 14152 9276 14216 9280
rect 14152 9220 14156 9276
rect 14156 9220 14212 9276
rect 14212 9220 14216 9276
rect 14152 9216 14216 9220
rect 14232 9276 14296 9280
rect 14232 9220 14236 9276
rect 14236 9220 14292 9276
rect 14292 9220 14296 9276
rect 14232 9216 14296 9220
rect 2652 8732 2716 8736
rect 2652 8676 2656 8732
rect 2656 8676 2712 8732
rect 2712 8676 2716 8732
rect 2652 8672 2716 8676
rect 2732 8732 2796 8736
rect 2732 8676 2736 8732
rect 2736 8676 2792 8732
rect 2792 8676 2796 8732
rect 2732 8672 2796 8676
rect 2812 8732 2876 8736
rect 2812 8676 2816 8732
rect 2816 8676 2872 8732
rect 2872 8676 2876 8732
rect 2812 8672 2876 8676
rect 2892 8732 2956 8736
rect 2892 8676 2896 8732
rect 2896 8676 2952 8732
rect 2952 8676 2956 8732
rect 2892 8672 2956 8676
rect 2972 8732 3036 8736
rect 2972 8676 2976 8732
rect 2976 8676 3032 8732
rect 3032 8676 3036 8732
rect 2972 8672 3036 8676
rect 8652 8732 8716 8736
rect 8652 8676 8656 8732
rect 8656 8676 8712 8732
rect 8712 8676 8716 8732
rect 8652 8672 8716 8676
rect 8732 8732 8796 8736
rect 8732 8676 8736 8732
rect 8736 8676 8792 8732
rect 8792 8676 8796 8732
rect 8732 8672 8796 8676
rect 8812 8732 8876 8736
rect 8812 8676 8816 8732
rect 8816 8676 8872 8732
rect 8872 8676 8876 8732
rect 8812 8672 8876 8676
rect 8892 8732 8956 8736
rect 8892 8676 8896 8732
rect 8896 8676 8952 8732
rect 8952 8676 8956 8732
rect 8892 8672 8956 8676
rect 8972 8732 9036 8736
rect 8972 8676 8976 8732
rect 8976 8676 9032 8732
rect 9032 8676 9036 8732
rect 8972 8672 9036 8676
rect 14652 8732 14716 8736
rect 14652 8676 14656 8732
rect 14656 8676 14712 8732
rect 14712 8676 14716 8732
rect 14652 8672 14716 8676
rect 14732 8732 14796 8736
rect 14732 8676 14736 8732
rect 14736 8676 14792 8732
rect 14792 8676 14796 8732
rect 14732 8672 14796 8676
rect 14812 8732 14876 8736
rect 14812 8676 14816 8732
rect 14816 8676 14872 8732
rect 14872 8676 14876 8732
rect 14812 8672 14876 8676
rect 14892 8732 14956 8736
rect 14892 8676 14896 8732
rect 14896 8676 14952 8732
rect 14952 8676 14956 8732
rect 14892 8672 14956 8676
rect 14972 8732 15036 8736
rect 14972 8676 14976 8732
rect 14976 8676 15032 8732
rect 15032 8676 15036 8732
rect 14972 8672 15036 8676
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 14152 8188 14216 8192
rect 14152 8132 14156 8188
rect 14156 8132 14212 8188
rect 14212 8132 14216 8188
rect 14152 8128 14216 8132
rect 14232 8188 14296 8192
rect 14232 8132 14236 8188
rect 14236 8132 14292 8188
rect 14292 8132 14296 8188
rect 14232 8128 14296 8132
rect 2652 7644 2716 7648
rect 2652 7588 2656 7644
rect 2656 7588 2712 7644
rect 2712 7588 2716 7644
rect 2652 7584 2716 7588
rect 2732 7644 2796 7648
rect 2732 7588 2736 7644
rect 2736 7588 2792 7644
rect 2792 7588 2796 7644
rect 2732 7584 2796 7588
rect 2812 7644 2876 7648
rect 2812 7588 2816 7644
rect 2816 7588 2872 7644
rect 2872 7588 2876 7644
rect 2812 7584 2876 7588
rect 2892 7644 2956 7648
rect 2892 7588 2896 7644
rect 2896 7588 2952 7644
rect 2952 7588 2956 7644
rect 2892 7584 2956 7588
rect 2972 7644 3036 7648
rect 2972 7588 2976 7644
rect 2976 7588 3032 7644
rect 3032 7588 3036 7644
rect 2972 7584 3036 7588
rect 8652 7644 8716 7648
rect 8652 7588 8656 7644
rect 8656 7588 8712 7644
rect 8712 7588 8716 7644
rect 8652 7584 8716 7588
rect 8732 7644 8796 7648
rect 8732 7588 8736 7644
rect 8736 7588 8792 7644
rect 8792 7588 8796 7644
rect 8732 7584 8796 7588
rect 8812 7644 8876 7648
rect 8812 7588 8816 7644
rect 8816 7588 8872 7644
rect 8872 7588 8876 7644
rect 8812 7584 8876 7588
rect 8892 7644 8956 7648
rect 8892 7588 8896 7644
rect 8896 7588 8952 7644
rect 8952 7588 8956 7644
rect 8892 7584 8956 7588
rect 8972 7644 9036 7648
rect 8972 7588 8976 7644
rect 8976 7588 9032 7644
rect 9032 7588 9036 7644
rect 8972 7584 9036 7588
rect 14652 7644 14716 7648
rect 14652 7588 14656 7644
rect 14656 7588 14712 7644
rect 14712 7588 14716 7644
rect 14652 7584 14716 7588
rect 14732 7644 14796 7648
rect 14732 7588 14736 7644
rect 14736 7588 14792 7644
rect 14792 7588 14796 7644
rect 14732 7584 14796 7588
rect 14812 7644 14876 7648
rect 14812 7588 14816 7644
rect 14816 7588 14872 7644
rect 14872 7588 14876 7644
rect 14812 7584 14876 7588
rect 14892 7644 14956 7648
rect 14892 7588 14896 7644
rect 14896 7588 14952 7644
rect 14952 7588 14956 7644
rect 14892 7584 14956 7588
rect 14972 7644 15036 7648
rect 14972 7588 14976 7644
rect 14976 7588 15032 7644
rect 15032 7588 15036 7644
rect 14972 7584 15036 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 14152 7100 14216 7104
rect 14152 7044 14156 7100
rect 14156 7044 14212 7100
rect 14212 7044 14216 7100
rect 14152 7040 14216 7044
rect 14232 7100 14296 7104
rect 14232 7044 14236 7100
rect 14236 7044 14292 7100
rect 14292 7044 14296 7100
rect 14232 7040 14296 7044
rect 2652 6556 2716 6560
rect 2652 6500 2656 6556
rect 2656 6500 2712 6556
rect 2712 6500 2716 6556
rect 2652 6496 2716 6500
rect 2732 6556 2796 6560
rect 2732 6500 2736 6556
rect 2736 6500 2792 6556
rect 2792 6500 2796 6556
rect 2732 6496 2796 6500
rect 2812 6556 2876 6560
rect 2812 6500 2816 6556
rect 2816 6500 2872 6556
rect 2872 6500 2876 6556
rect 2812 6496 2876 6500
rect 2892 6556 2956 6560
rect 2892 6500 2896 6556
rect 2896 6500 2952 6556
rect 2952 6500 2956 6556
rect 2892 6496 2956 6500
rect 2972 6556 3036 6560
rect 2972 6500 2976 6556
rect 2976 6500 3032 6556
rect 3032 6500 3036 6556
rect 2972 6496 3036 6500
rect 8652 6556 8716 6560
rect 8652 6500 8656 6556
rect 8656 6500 8712 6556
rect 8712 6500 8716 6556
rect 8652 6496 8716 6500
rect 8732 6556 8796 6560
rect 8732 6500 8736 6556
rect 8736 6500 8792 6556
rect 8792 6500 8796 6556
rect 8732 6496 8796 6500
rect 8812 6556 8876 6560
rect 8812 6500 8816 6556
rect 8816 6500 8872 6556
rect 8872 6500 8876 6556
rect 8812 6496 8876 6500
rect 8892 6556 8956 6560
rect 8892 6500 8896 6556
rect 8896 6500 8952 6556
rect 8952 6500 8956 6556
rect 8892 6496 8956 6500
rect 8972 6556 9036 6560
rect 8972 6500 8976 6556
rect 8976 6500 9032 6556
rect 9032 6500 9036 6556
rect 8972 6496 9036 6500
rect 14652 6556 14716 6560
rect 14652 6500 14656 6556
rect 14656 6500 14712 6556
rect 14712 6500 14716 6556
rect 14652 6496 14716 6500
rect 14732 6556 14796 6560
rect 14732 6500 14736 6556
rect 14736 6500 14792 6556
rect 14792 6500 14796 6556
rect 14732 6496 14796 6500
rect 14812 6556 14876 6560
rect 14812 6500 14816 6556
rect 14816 6500 14872 6556
rect 14872 6500 14876 6556
rect 14812 6496 14876 6500
rect 14892 6556 14956 6560
rect 14892 6500 14896 6556
rect 14896 6500 14952 6556
rect 14952 6500 14956 6556
rect 14892 6496 14956 6500
rect 14972 6556 15036 6560
rect 14972 6500 14976 6556
rect 14976 6500 15032 6556
rect 15032 6500 15036 6556
rect 14972 6496 15036 6500
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 14152 6012 14216 6016
rect 14152 5956 14156 6012
rect 14156 5956 14212 6012
rect 14212 5956 14216 6012
rect 14152 5952 14216 5956
rect 14232 6012 14296 6016
rect 14232 5956 14236 6012
rect 14236 5956 14292 6012
rect 14292 5956 14296 6012
rect 14232 5952 14296 5956
rect 16620 5808 16684 5812
rect 16620 5752 16634 5808
rect 16634 5752 16684 5808
rect 16620 5748 16684 5752
rect 2652 5468 2716 5472
rect 2652 5412 2656 5468
rect 2656 5412 2712 5468
rect 2712 5412 2716 5468
rect 2652 5408 2716 5412
rect 2732 5468 2796 5472
rect 2732 5412 2736 5468
rect 2736 5412 2792 5468
rect 2792 5412 2796 5468
rect 2732 5408 2796 5412
rect 2812 5468 2876 5472
rect 2812 5412 2816 5468
rect 2816 5412 2872 5468
rect 2872 5412 2876 5468
rect 2812 5408 2876 5412
rect 2892 5468 2956 5472
rect 2892 5412 2896 5468
rect 2896 5412 2952 5468
rect 2952 5412 2956 5468
rect 2892 5408 2956 5412
rect 2972 5468 3036 5472
rect 2972 5412 2976 5468
rect 2976 5412 3032 5468
rect 3032 5412 3036 5468
rect 2972 5408 3036 5412
rect 8652 5468 8716 5472
rect 8652 5412 8656 5468
rect 8656 5412 8712 5468
rect 8712 5412 8716 5468
rect 8652 5408 8716 5412
rect 8732 5468 8796 5472
rect 8732 5412 8736 5468
rect 8736 5412 8792 5468
rect 8792 5412 8796 5468
rect 8732 5408 8796 5412
rect 8812 5468 8876 5472
rect 8812 5412 8816 5468
rect 8816 5412 8872 5468
rect 8872 5412 8876 5468
rect 8812 5408 8876 5412
rect 8892 5468 8956 5472
rect 8892 5412 8896 5468
rect 8896 5412 8952 5468
rect 8952 5412 8956 5468
rect 8892 5408 8956 5412
rect 8972 5468 9036 5472
rect 8972 5412 8976 5468
rect 8976 5412 9032 5468
rect 9032 5412 9036 5468
rect 8972 5408 9036 5412
rect 14652 5468 14716 5472
rect 14652 5412 14656 5468
rect 14656 5412 14712 5468
rect 14712 5412 14716 5468
rect 14652 5408 14716 5412
rect 14732 5468 14796 5472
rect 14732 5412 14736 5468
rect 14736 5412 14792 5468
rect 14792 5412 14796 5468
rect 14732 5408 14796 5412
rect 14812 5468 14876 5472
rect 14812 5412 14816 5468
rect 14816 5412 14872 5468
rect 14872 5412 14876 5468
rect 14812 5408 14876 5412
rect 14892 5468 14956 5472
rect 14892 5412 14896 5468
rect 14896 5412 14952 5468
rect 14952 5412 14956 5468
rect 14892 5408 14956 5412
rect 14972 5468 15036 5472
rect 14972 5412 14976 5468
rect 14976 5412 15032 5468
rect 15032 5412 15036 5468
rect 14972 5408 15036 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 14152 4924 14216 4928
rect 14152 4868 14156 4924
rect 14156 4868 14212 4924
rect 14212 4868 14216 4924
rect 14152 4864 14216 4868
rect 14232 4924 14296 4928
rect 14232 4868 14236 4924
rect 14236 4868 14292 4924
rect 14292 4868 14296 4924
rect 14232 4864 14296 4868
rect 2652 4380 2716 4384
rect 2652 4324 2656 4380
rect 2656 4324 2712 4380
rect 2712 4324 2716 4380
rect 2652 4320 2716 4324
rect 2732 4380 2796 4384
rect 2732 4324 2736 4380
rect 2736 4324 2792 4380
rect 2792 4324 2796 4380
rect 2732 4320 2796 4324
rect 2812 4380 2876 4384
rect 2812 4324 2816 4380
rect 2816 4324 2872 4380
rect 2872 4324 2876 4380
rect 2812 4320 2876 4324
rect 2892 4380 2956 4384
rect 2892 4324 2896 4380
rect 2896 4324 2952 4380
rect 2952 4324 2956 4380
rect 2892 4320 2956 4324
rect 2972 4380 3036 4384
rect 2972 4324 2976 4380
rect 2976 4324 3032 4380
rect 3032 4324 3036 4380
rect 2972 4320 3036 4324
rect 8652 4380 8716 4384
rect 8652 4324 8656 4380
rect 8656 4324 8712 4380
rect 8712 4324 8716 4380
rect 8652 4320 8716 4324
rect 8732 4380 8796 4384
rect 8732 4324 8736 4380
rect 8736 4324 8792 4380
rect 8792 4324 8796 4380
rect 8732 4320 8796 4324
rect 8812 4380 8876 4384
rect 8812 4324 8816 4380
rect 8816 4324 8872 4380
rect 8872 4324 8876 4380
rect 8812 4320 8876 4324
rect 8892 4380 8956 4384
rect 8892 4324 8896 4380
rect 8896 4324 8952 4380
rect 8952 4324 8956 4380
rect 8892 4320 8956 4324
rect 8972 4380 9036 4384
rect 8972 4324 8976 4380
rect 8976 4324 9032 4380
rect 9032 4324 9036 4380
rect 8972 4320 9036 4324
rect 14652 4380 14716 4384
rect 14652 4324 14656 4380
rect 14656 4324 14712 4380
rect 14712 4324 14716 4380
rect 14652 4320 14716 4324
rect 14732 4380 14796 4384
rect 14732 4324 14736 4380
rect 14736 4324 14792 4380
rect 14792 4324 14796 4380
rect 14732 4320 14796 4324
rect 14812 4380 14876 4384
rect 14812 4324 14816 4380
rect 14816 4324 14872 4380
rect 14872 4324 14876 4380
rect 14812 4320 14876 4324
rect 14892 4380 14956 4384
rect 14892 4324 14896 4380
rect 14896 4324 14952 4380
rect 14952 4324 14956 4380
rect 14892 4320 14956 4324
rect 14972 4380 15036 4384
rect 14972 4324 14976 4380
rect 14976 4324 15032 4380
rect 15032 4324 15036 4380
rect 14972 4320 15036 4324
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 14152 3836 14216 3840
rect 14152 3780 14156 3836
rect 14156 3780 14212 3836
rect 14212 3780 14216 3836
rect 14152 3776 14216 3780
rect 14232 3836 14296 3840
rect 14232 3780 14236 3836
rect 14236 3780 14292 3836
rect 14292 3780 14296 3836
rect 14232 3776 14296 3780
rect 2652 3292 2716 3296
rect 2652 3236 2656 3292
rect 2656 3236 2712 3292
rect 2712 3236 2716 3292
rect 2652 3232 2716 3236
rect 2732 3292 2796 3296
rect 2732 3236 2736 3292
rect 2736 3236 2792 3292
rect 2792 3236 2796 3292
rect 2732 3232 2796 3236
rect 2812 3292 2876 3296
rect 2812 3236 2816 3292
rect 2816 3236 2872 3292
rect 2872 3236 2876 3292
rect 2812 3232 2876 3236
rect 2892 3292 2956 3296
rect 2892 3236 2896 3292
rect 2896 3236 2952 3292
rect 2952 3236 2956 3292
rect 2892 3232 2956 3236
rect 2972 3292 3036 3296
rect 2972 3236 2976 3292
rect 2976 3236 3032 3292
rect 3032 3236 3036 3292
rect 2972 3232 3036 3236
rect 8652 3292 8716 3296
rect 8652 3236 8656 3292
rect 8656 3236 8712 3292
rect 8712 3236 8716 3292
rect 8652 3232 8716 3236
rect 8732 3292 8796 3296
rect 8732 3236 8736 3292
rect 8736 3236 8792 3292
rect 8792 3236 8796 3292
rect 8732 3232 8796 3236
rect 8812 3292 8876 3296
rect 8812 3236 8816 3292
rect 8816 3236 8872 3292
rect 8872 3236 8876 3292
rect 8812 3232 8876 3236
rect 8892 3292 8956 3296
rect 8892 3236 8896 3292
rect 8896 3236 8952 3292
rect 8952 3236 8956 3292
rect 8892 3232 8956 3236
rect 8972 3292 9036 3296
rect 8972 3236 8976 3292
rect 8976 3236 9032 3292
rect 9032 3236 9036 3292
rect 8972 3232 9036 3236
rect 14652 3292 14716 3296
rect 14652 3236 14656 3292
rect 14656 3236 14712 3292
rect 14712 3236 14716 3292
rect 14652 3232 14716 3236
rect 14732 3292 14796 3296
rect 14732 3236 14736 3292
rect 14736 3236 14792 3292
rect 14792 3236 14796 3292
rect 14732 3232 14796 3236
rect 14812 3292 14876 3296
rect 14812 3236 14816 3292
rect 14816 3236 14872 3292
rect 14872 3236 14876 3292
rect 14812 3232 14876 3236
rect 14892 3292 14956 3296
rect 14892 3236 14896 3292
rect 14896 3236 14952 3292
rect 14952 3236 14956 3292
rect 14892 3232 14956 3236
rect 14972 3292 15036 3296
rect 14972 3236 14976 3292
rect 14976 3236 15032 3292
rect 15032 3236 15036 3292
rect 14972 3232 15036 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 14152 2748 14216 2752
rect 14152 2692 14156 2748
rect 14156 2692 14212 2748
rect 14212 2692 14216 2748
rect 14152 2688 14216 2692
rect 14232 2748 14296 2752
rect 14232 2692 14236 2748
rect 14236 2692 14292 2748
rect 14292 2692 14296 2748
rect 14232 2688 14296 2692
rect 2652 2204 2716 2208
rect 2652 2148 2656 2204
rect 2656 2148 2712 2204
rect 2712 2148 2716 2204
rect 2652 2144 2716 2148
rect 2732 2204 2796 2208
rect 2732 2148 2736 2204
rect 2736 2148 2792 2204
rect 2792 2148 2796 2204
rect 2732 2144 2796 2148
rect 2812 2204 2876 2208
rect 2812 2148 2816 2204
rect 2816 2148 2872 2204
rect 2872 2148 2876 2204
rect 2812 2144 2876 2148
rect 2892 2204 2956 2208
rect 2892 2148 2896 2204
rect 2896 2148 2952 2204
rect 2952 2148 2956 2204
rect 2892 2144 2956 2148
rect 2972 2204 3036 2208
rect 2972 2148 2976 2204
rect 2976 2148 3032 2204
rect 3032 2148 3036 2204
rect 2972 2144 3036 2148
rect 8652 2204 8716 2208
rect 8652 2148 8656 2204
rect 8656 2148 8712 2204
rect 8712 2148 8716 2204
rect 8652 2144 8716 2148
rect 8732 2204 8796 2208
rect 8732 2148 8736 2204
rect 8736 2148 8792 2204
rect 8792 2148 8796 2204
rect 8732 2144 8796 2148
rect 8812 2204 8876 2208
rect 8812 2148 8816 2204
rect 8816 2148 8872 2204
rect 8872 2148 8876 2204
rect 8812 2144 8876 2148
rect 8892 2204 8956 2208
rect 8892 2148 8896 2204
rect 8896 2148 8952 2204
rect 8952 2148 8956 2204
rect 8892 2144 8956 2148
rect 8972 2204 9036 2208
rect 8972 2148 8976 2204
rect 8976 2148 9032 2204
rect 9032 2148 9036 2204
rect 8972 2144 9036 2148
rect 14652 2204 14716 2208
rect 14652 2148 14656 2204
rect 14656 2148 14712 2204
rect 14712 2148 14716 2204
rect 14652 2144 14716 2148
rect 14732 2204 14796 2208
rect 14732 2148 14736 2204
rect 14736 2148 14792 2204
rect 14792 2148 14796 2204
rect 14732 2144 14796 2148
rect 14812 2204 14876 2208
rect 14812 2148 14816 2204
rect 14816 2148 14872 2204
rect 14872 2148 14876 2204
rect 14812 2144 14876 2148
rect 14892 2204 14956 2208
rect 14892 2148 14896 2204
rect 14896 2148 14952 2204
rect 14952 2148 14956 2204
rect 14892 2144 14956 2148
rect 14972 2204 15036 2208
rect 14972 2148 14976 2204
rect 14976 2148 15032 2204
rect 15032 2148 15036 2204
rect 14972 2144 15036 2148
<< metal4 >>
rect 1904 19072 2304 19088
rect 1904 19008 1912 19072
rect 1976 19008 1992 19072
rect 2056 19008 2072 19072
rect 2136 19008 2152 19072
rect 2216 19008 2232 19072
rect 2296 19008 2304 19072
rect 1904 17984 2304 19008
rect 1904 17920 1912 17984
rect 1976 17920 1992 17984
rect 2056 17920 2072 17984
rect 2136 17920 2152 17984
rect 2216 17920 2232 17984
rect 2296 17920 2304 17984
rect 1904 16896 2304 17920
rect 1904 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2304 16896
rect 1904 15808 2304 16832
rect 1904 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2304 15808
rect 1904 15294 2304 15744
rect 1904 15058 1986 15294
rect 2222 15058 2304 15294
rect 1904 14720 2304 15058
rect 1904 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2304 14720
rect 1904 13632 2304 14656
rect 1904 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2304 13632
rect 1904 12544 2304 13568
rect 1904 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2304 12544
rect 1904 11456 2304 12480
rect 1904 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2304 11456
rect 1904 10368 2304 11392
rect 1904 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2304 10368
rect 1904 9294 2304 10304
rect 1904 9280 1986 9294
rect 2222 9280 2304 9294
rect 1904 9216 1912 9280
rect 1976 9216 1986 9280
rect 2222 9216 2232 9280
rect 2296 9216 2304 9280
rect 1904 9058 1986 9216
rect 2222 9058 2304 9216
rect 1904 8192 2304 9058
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 3294 2304 3776
rect 1904 3058 1986 3294
rect 2222 3058 2304 3294
rect 1904 2752 2304 3058
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 2128 2304 2688
rect 2644 18528 3044 19088
rect 2644 18464 2652 18528
rect 2716 18464 2732 18528
rect 2796 18464 2812 18528
rect 2876 18464 2892 18528
rect 2956 18464 2972 18528
rect 3036 18464 3044 18528
rect 2644 17440 3044 18464
rect 2644 17376 2652 17440
rect 2716 17376 2732 17440
rect 2796 17376 2812 17440
rect 2876 17376 2892 17440
rect 2956 17376 2972 17440
rect 3036 17376 3044 17440
rect 2644 16352 3044 17376
rect 2644 16288 2652 16352
rect 2716 16288 2732 16352
rect 2796 16288 2812 16352
rect 2876 16288 2892 16352
rect 2956 16288 2972 16352
rect 3036 16288 3044 16352
rect 2644 16034 3044 16288
rect 2644 15798 2726 16034
rect 2962 15798 3044 16034
rect 2644 15264 3044 15798
rect 2644 15200 2652 15264
rect 2716 15200 2732 15264
rect 2796 15200 2812 15264
rect 2876 15200 2892 15264
rect 2956 15200 2972 15264
rect 3036 15200 3044 15264
rect 2644 14176 3044 15200
rect 2644 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3044 14176
rect 2644 13088 3044 14112
rect 2644 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3044 13088
rect 2644 12000 3044 13024
rect 2644 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3044 12000
rect 2644 10912 3044 11936
rect 2644 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3044 10912
rect 2644 10034 3044 10848
rect 2644 9824 2726 10034
rect 2962 9824 3044 10034
rect 2644 9760 2652 9824
rect 2716 9798 2726 9824
rect 2962 9798 2972 9824
rect 2716 9760 2732 9798
rect 2796 9760 2812 9798
rect 2876 9760 2892 9798
rect 2956 9760 2972 9798
rect 3036 9760 3044 9824
rect 2644 8736 3044 9760
rect 2644 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3044 8736
rect 2644 7648 3044 8672
rect 2644 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3044 7648
rect 2644 6560 3044 7584
rect 2644 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3044 6560
rect 2644 5472 3044 6496
rect 2644 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3044 5472
rect 2644 4384 3044 5408
rect 2644 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3044 4384
rect 2644 4034 3044 4320
rect 2644 3798 2726 4034
rect 2962 3798 3044 4034
rect 2644 3296 3044 3798
rect 2644 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3044 3296
rect 2644 2208 3044 3232
rect 2644 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3044 2208
rect 2644 2128 3044 2144
rect 7904 19072 8304 19088
rect 7904 19008 7912 19072
rect 7976 19008 7992 19072
rect 8056 19008 8072 19072
rect 8136 19008 8152 19072
rect 8216 19008 8232 19072
rect 8296 19008 8304 19072
rect 7904 17984 8304 19008
rect 7904 17920 7912 17984
rect 7976 17920 7992 17984
rect 8056 17920 8072 17984
rect 8136 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8304 17984
rect 7904 16896 8304 17920
rect 7904 16832 7912 16896
rect 7976 16832 7992 16896
rect 8056 16832 8072 16896
rect 8136 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8304 16896
rect 7904 15808 8304 16832
rect 7904 15744 7912 15808
rect 7976 15744 7992 15808
rect 8056 15744 8072 15808
rect 8136 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8304 15808
rect 7904 15294 8304 15744
rect 7904 15058 7986 15294
rect 8222 15058 8304 15294
rect 7904 14720 8304 15058
rect 7904 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8304 14720
rect 7904 13632 8304 14656
rect 7904 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8304 13632
rect 7904 12544 8304 13568
rect 7904 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8304 12544
rect 7904 11456 8304 12480
rect 7904 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8304 11456
rect 7904 10368 8304 11392
rect 7904 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8304 10368
rect 7904 9294 8304 10304
rect 7904 9280 7986 9294
rect 8222 9280 8304 9294
rect 7904 9216 7912 9280
rect 7976 9216 7986 9280
rect 8222 9216 8232 9280
rect 8296 9216 8304 9280
rect 7904 9058 7986 9216
rect 8222 9058 8304 9216
rect 7904 8192 8304 9058
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 7904 7104 8304 8128
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 7904 3840 8304 4864
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 3294 8304 3776
rect 7904 3058 7986 3294
rect 8222 3058 8304 3294
rect 7904 2752 8304 3058
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 2128 8304 2688
rect 8644 18528 9044 19088
rect 8644 18464 8652 18528
rect 8716 18464 8732 18528
rect 8796 18464 8812 18528
rect 8876 18464 8892 18528
rect 8956 18464 8972 18528
rect 9036 18464 9044 18528
rect 8644 17440 9044 18464
rect 8644 17376 8652 17440
rect 8716 17376 8732 17440
rect 8796 17376 8812 17440
rect 8876 17376 8892 17440
rect 8956 17376 8972 17440
rect 9036 17376 9044 17440
rect 8644 16352 9044 17376
rect 8644 16288 8652 16352
rect 8716 16288 8732 16352
rect 8796 16288 8812 16352
rect 8876 16288 8892 16352
rect 8956 16288 8972 16352
rect 9036 16288 9044 16352
rect 8644 16034 9044 16288
rect 8644 15798 8726 16034
rect 8962 15798 9044 16034
rect 8644 15264 9044 15798
rect 8644 15200 8652 15264
rect 8716 15200 8732 15264
rect 8796 15200 8812 15264
rect 8876 15200 8892 15264
rect 8956 15200 8972 15264
rect 9036 15200 9044 15264
rect 8644 14176 9044 15200
rect 8644 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9044 14176
rect 8644 13088 9044 14112
rect 8644 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9044 13088
rect 8644 12000 9044 13024
rect 8644 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9044 12000
rect 8644 10912 9044 11936
rect 8644 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9044 10912
rect 8644 10034 9044 10848
rect 8644 9824 8726 10034
rect 8962 9824 9044 10034
rect 8644 9760 8652 9824
rect 8716 9798 8726 9824
rect 8962 9798 8972 9824
rect 8716 9760 8732 9798
rect 8796 9760 8812 9798
rect 8876 9760 8892 9798
rect 8956 9760 8972 9798
rect 9036 9760 9044 9824
rect 8644 8736 9044 9760
rect 8644 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9044 8736
rect 8644 7648 9044 8672
rect 8644 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9044 7648
rect 8644 6560 9044 7584
rect 8644 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9044 6560
rect 8644 5472 9044 6496
rect 8644 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9044 5472
rect 8644 4384 9044 5408
rect 8644 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9044 4384
rect 8644 4034 9044 4320
rect 8644 3798 8726 4034
rect 8962 3798 9044 4034
rect 8644 3296 9044 3798
rect 8644 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9044 3296
rect 8644 2208 9044 3232
rect 8644 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9044 2208
rect 8644 2128 9044 2144
rect 13904 19072 14304 19088
rect 13904 19008 13912 19072
rect 13976 19008 13992 19072
rect 14056 19008 14072 19072
rect 14136 19008 14152 19072
rect 14216 19008 14232 19072
rect 14296 19008 14304 19072
rect 13904 17984 14304 19008
rect 13904 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14152 17984
rect 14216 17920 14232 17984
rect 14296 17920 14304 17984
rect 13904 16896 14304 17920
rect 13904 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14152 16896
rect 14216 16832 14232 16896
rect 14296 16832 14304 16896
rect 13904 15808 14304 16832
rect 13904 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14152 15808
rect 14216 15744 14232 15808
rect 14296 15744 14304 15808
rect 13904 15294 14304 15744
rect 13904 15058 13986 15294
rect 14222 15058 14304 15294
rect 13904 14720 14304 15058
rect 13904 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14304 14720
rect 13904 13632 14304 14656
rect 13904 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14304 13632
rect 13904 12544 14304 13568
rect 13904 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14304 12544
rect 13904 11456 14304 12480
rect 13904 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14304 11456
rect 13904 10368 14304 11392
rect 13904 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14304 10368
rect 13904 9294 14304 10304
rect 13904 9280 13986 9294
rect 14222 9280 14304 9294
rect 13904 9216 13912 9280
rect 13976 9216 13986 9280
rect 14222 9216 14232 9280
rect 14296 9216 14304 9280
rect 13904 9058 13986 9216
rect 14222 9058 14304 9216
rect 13904 8192 14304 9058
rect 13904 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14304 8192
rect 13904 7104 14304 8128
rect 13904 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14304 7104
rect 13904 6016 14304 7040
rect 13904 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14304 6016
rect 13904 4928 14304 5952
rect 13904 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14304 4928
rect 13904 3840 14304 4864
rect 13904 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14304 3840
rect 13904 3294 14304 3776
rect 13904 3058 13986 3294
rect 14222 3058 14304 3294
rect 13904 2752 14304 3058
rect 13904 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14304 2752
rect 13904 2128 14304 2688
rect 14644 18528 15044 19088
rect 14644 18464 14652 18528
rect 14716 18464 14732 18528
rect 14796 18464 14812 18528
rect 14876 18464 14892 18528
rect 14956 18464 14972 18528
rect 15036 18464 15044 18528
rect 14644 17440 15044 18464
rect 16619 18052 16685 18053
rect 16619 17988 16620 18052
rect 16684 17988 16685 18052
rect 16619 17987 16685 17988
rect 14644 17376 14652 17440
rect 14716 17376 14732 17440
rect 14796 17376 14812 17440
rect 14876 17376 14892 17440
rect 14956 17376 14972 17440
rect 15036 17376 15044 17440
rect 14644 16352 15044 17376
rect 14644 16288 14652 16352
rect 14716 16288 14732 16352
rect 14796 16288 14812 16352
rect 14876 16288 14892 16352
rect 14956 16288 14972 16352
rect 15036 16288 15044 16352
rect 14644 16034 15044 16288
rect 14644 15798 14726 16034
rect 14962 15798 15044 16034
rect 14644 15264 15044 15798
rect 14644 15200 14652 15264
rect 14716 15200 14732 15264
rect 14796 15200 14812 15264
rect 14876 15200 14892 15264
rect 14956 15200 14972 15264
rect 15036 15200 15044 15264
rect 14644 14176 15044 15200
rect 14644 14112 14652 14176
rect 14716 14112 14732 14176
rect 14796 14112 14812 14176
rect 14876 14112 14892 14176
rect 14956 14112 14972 14176
rect 15036 14112 15044 14176
rect 14644 13088 15044 14112
rect 14644 13024 14652 13088
rect 14716 13024 14732 13088
rect 14796 13024 14812 13088
rect 14876 13024 14892 13088
rect 14956 13024 14972 13088
rect 15036 13024 15044 13088
rect 14644 12000 15044 13024
rect 14644 11936 14652 12000
rect 14716 11936 14732 12000
rect 14796 11936 14812 12000
rect 14876 11936 14892 12000
rect 14956 11936 14972 12000
rect 15036 11936 15044 12000
rect 14644 10912 15044 11936
rect 14644 10848 14652 10912
rect 14716 10848 14732 10912
rect 14796 10848 14812 10912
rect 14876 10848 14892 10912
rect 14956 10848 14972 10912
rect 15036 10848 15044 10912
rect 14644 10034 15044 10848
rect 14644 9824 14726 10034
rect 14962 9824 15044 10034
rect 14644 9760 14652 9824
rect 14716 9798 14726 9824
rect 14962 9798 14972 9824
rect 14716 9760 14732 9798
rect 14796 9760 14812 9798
rect 14876 9760 14892 9798
rect 14956 9760 14972 9798
rect 15036 9760 15044 9824
rect 14644 8736 15044 9760
rect 14644 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15044 8736
rect 14644 7648 15044 8672
rect 14644 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15044 7648
rect 14644 6560 15044 7584
rect 14644 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15044 6560
rect 14644 5472 15044 6496
rect 16622 5813 16682 17987
rect 16619 5812 16685 5813
rect 16619 5748 16620 5812
rect 16684 5748 16685 5812
rect 16619 5747 16685 5748
rect 14644 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15044 5472
rect 14644 4384 15044 5408
rect 14644 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15044 4384
rect 14644 4034 15044 4320
rect 14644 3798 14726 4034
rect 14962 3798 15044 4034
rect 14644 3296 15044 3798
rect 14644 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15044 3296
rect 14644 2208 15044 3232
rect 14644 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15044 2208
rect 14644 2128 15044 2144
<< via4 >>
rect 1986 15058 2222 15294
rect 1986 9280 2222 9294
rect 1986 9216 1992 9280
rect 1992 9216 2056 9280
rect 2056 9216 2072 9280
rect 2072 9216 2136 9280
rect 2136 9216 2152 9280
rect 2152 9216 2216 9280
rect 2216 9216 2222 9280
rect 1986 9058 2222 9216
rect 1986 3058 2222 3294
rect 2726 15798 2962 16034
rect 2726 9824 2962 10034
rect 2726 9798 2732 9824
rect 2732 9798 2796 9824
rect 2796 9798 2812 9824
rect 2812 9798 2876 9824
rect 2876 9798 2892 9824
rect 2892 9798 2956 9824
rect 2956 9798 2962 9824
rect 2726 3798 2962 4034
rect 7986 15058 8222 15294
rect 7986 9280 8222 9294
rect 7986 9216 7992 9280
rect 7992 9216 8056 9280
rect 8056 9216 8072 9280
rect 8072 9216 8136 9280
rect 8136 9216 8152 9280
rect 8152 9216 8216 9280
rect 8216 9216 8222 9280
rect 7986 9058 8222 9216
rect 7986 3058 8222 3294
rect 8726 15798 8962 16034
rect 8726 9824 8962 10034
rect 8726 9798 8732 9824
rect 8732 9798 8796 9824
rect 8796 9798 8812 9824
rect 8812 9798 8876 9824
rect 8876 9798 8892 9824
rect 8892 9798 8956 9824
rect 8956 9798 8962 9824
rect 8726 3798 8962 4034
rect 13986 15058 14222 15294
rect 13986 9280 14222 9294
rect 13986 9216 13992 9280
rect 13992 9216 14056 9280
rect 14056 9216 14072 9280
rect 14072 9216 14136 9280
rect 14136 9216 14152 9280
rect 14152 9216 14216 9280
rect 14216 9216 14222 9280
rect 13986 9058 14222 9216
rect 13986 3058 14222 3294
rect 14726 15798 14962 16034
rect 14726 9824 14962 10034
rect 14726 9798 14732 9824
rect 14732 9798 14796 9824
rect 14796 9798 14812 9824
rect 14812 9798 14876 9824
rect 14876 9798 14892 9824
rect 14892 9798 14956 9824
rect 14956 9798 14962 9824
rect 14726 3798 14962 4034
<< metal5 >>
rect 1056 16034 18264 16116
rect 1056 15798 2726 16034
rect 2962 15798 8726 16034
rect 8962 15798 14726 16034
rect 14962 15798 18264 16034
rect 1056 15716 18264 15798
rect 1056 15294 18264 15376
rect 1056 15058 1986 15294
rect 2222 15058 7986 15294
rect 8222 15058 13986 15294
rect 14222 15058 18264 15294
rect 1056 14976 18264 15058
rect 1056 10034 18264 10116
rect 1056 9798 2726 10034
rect 2962 9798 8726 10034
rect 8962 9798 14726 10034
rect 14962 9798 18264 10034
rect 1056 9716 18264 9798
rect 1056 9294 18264 9376
rect 1056 9058 1986 9294
rect 2222 9058 7986 9294
rect 8222 9058 13986 9294
rect 14222 9058 18264 9294
rect 1056 8976 18264 9058
rect 1056 4034 18264 4116
rect 1056 3798 2726 4034
rect 2962 3798 8726 4034
rect 8962 3798 14726 4034
rect 14962 3798 18264 4034
rect 1056 3716 18264 3798
rect 1056 3294 18264 3376
rect 1056 3058 1986 3294
rect 2222 3058 7986 3294
rect 8222 3058 13986 3294
rect 14222 3058 18264 3294
rect 1056 2976 18264 3058
use sky130_fd_sc_hd__clkbuf_4  _102_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _103_
timestamp 0
transform -1 0 13892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _104_
timestamp 0
transform -1 0 12880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _105_
timestamp 0
transform 1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _106_
timestamp 0
transform 1 0 12788 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 0
transform -1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _108_
timestamp 0
transform -1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _109_
timestamp 0
transform 1 0 7636 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _110_
timestamp 0
transform -1 0 8004 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _111_
timestamp 0
transform 1 0 12972 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _112_
timestamp 0
transform 1 0 6164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _113_
timestamp 0
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _114_
timestamp 0
transform -1 0 12972 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _115_
timestamp 0
transform -1 0 11776 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _116_
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _117_
timestamp 0
transform -1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _118_
timestamp 0
transform 1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _119_
timestamp 0
transform 1 0 1472 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _120_
timestamp 0
transform -1 0 15548 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _121_
timestamp 0
transform 1 0 15548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _122_
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _123_
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _124_
timestamp 0
transform 1 0 4784 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _125_
timestamp 0
transform -1 0 5704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _126_
timestamp 0
transform -1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _127_
timestamp 0
transform -1 0 4968 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _128_
timestamp 0
transform 1 0 15088 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _129_
timestamp 0
transform -1 0 16008 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _130_
timestamp 0
transform -1 0 14904 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _131_
timestamp 0
transform -1 0 14812 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _132_
timestamp 0
transform -1 0 3312 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _133_
timestamp 0
transform -1 0 2760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _134_
timestamp 0
transform -1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _135_
timestamp 0
transform 1 0 3128 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _136_
timestamp 0
transform 1 0 15088 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _137_
timestamp 0
transform -1 0 16008 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _138_
timestamp 0
transform -1 0 14904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _139_
timestamp 0
transform 1 0 14168 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _140_
timestamp 0
transform 1 0 3220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _141_
timestamp 0
transform -1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _142_
timestamp 0
transform 1 0 3128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _143_
timestamp 0
transform 1 0 2576 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _144_
timestamp 0
transform 1 0 6716 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _145_
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _146_
timestamp 0
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _147_
timestamp 0
transform -1 0 15272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _148_
timestamp 0
transform -1 0 14720 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _149_
timestamp 0
transform -1 0 16560 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _150_
timestamp 0
transform -1 0 16836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _151_
timestamp 0
transform 1 0 16744 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _152_
timestamp 0
transform -1 0 17480 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _153_
timestamp 0
transform 1 0 2944 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _154_
timestamp 0
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _155_
timestamp 0
transform -1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _156_
timestamp 0
transform -1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _157_
timestamp 0
transform -1 0 2668 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _158_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _159_
timestamp 0
transform -1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _160_
timestamp 0
transform 1 0 3496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _161_
timestamp 0
transform -1 0 4232 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _162_
timestamp 0
transform -1 0 5152 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _163_
timestamp 0
transform -1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _164_
timestamp 0
transform -1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _165_
timestamp 0
transform 1 0 4048 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _166_
timestamp 0
transform -1 0 12236 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _167_
timestamp 0
transform -1 0 11408 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _168_
timestamp 0
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _169_
timestamp 0
transform -1 0 13340 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _170_
timestamp 0
transform 1 0 10764 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _171_
timestamp 0
transform -1 0 10304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _172_
timestamp 0
transform 1 0 10580 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _173_
timestamp 0
transform -1 0 10580 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _174_
timestamp 0
transform 1 0 7176 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _175_
timestamp 0
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _176_
timestamp 0
transform -1 0 6992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _177_
timestamp 0
transform 1 0 5060 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _178_
timestamp 0
transform -1 0 5612 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _179_
timestamp 0
transform -1 0 5152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _180_
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _181_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _182_
timestamp 0
transform -1 0 11224 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _183_
timestamp 0
transform -1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _184_
timestamp 0
transform -1 0 11500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _185_
timestamp 0
transform -1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _186_
timestamp 0
transform 1 0 17020 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 0
transform -1 0 17756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _188_
timestamp 0
transform 1 0 16744 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _189_
timestamp 0
transform 1 0 17112 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _190_
timestamp 0
transform -1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _191_
timestamp 0
transform -1 0 10580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _192_
timestamp 0
transform -1 0 11500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _193_
timestamp 0
transform 1 0 10212 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _194_
timestamp 0
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _195_
timestamp 0
transform -1 0 5520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _196_
timestamp 0
transform 1 0 5612 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _197_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _198_
timestamp 0
transform -1 0 10212 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _199_
timestamp 0
transform -1 0 17020 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _200_
timestamp 0
transform -1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _201_
timestamp 0
transform -1 0 8924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _202_
timestamp 0
transform -1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _203_
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _204_
timestamp 0
transform -1 0 12696 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _205_
timestamp 0
transform -1 0 12972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _206_
timestamp 0
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _207_
timestamp 0
transform -1 0 12788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _208_
timestamp 0
transform -1 0 7636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _209_
timestamp 0
transform -1 0 12696 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _210_
timestamp 0
transform -1 0 2392 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _211_
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _212_
timestamp 0
transform -1 0 5152 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _213_
timestamp 0
transform -1 0 15088 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _214_
timestamp 0
transform -1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 0
transform -1 0 15088 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _216_
timestamp 0
transform -1 0 3128 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _217_
timestamp 0
transform -1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _218_
timestamp 0
transform -1 0 16468 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _219_
timestamp 0
transform -1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _220_
timestamp 0
transform -1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _221_
timestamp 0
transform -1 0 4876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _222_
timestamp 0
transform -1 0 12696 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _223_
timestamp 0
transform -1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _224_
timestamp 0
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _225_
timestamp 0
transform -1 0 5796 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _226_
timestamp 0
transform -1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _227_
timestamp 0
transform -1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _228_
timestamp 0
transform -1 0 5796 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _229_
timestamp 0
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _230_
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _231_
timestamp 0
transform 1 0 10212 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 0
transform -1 0 11132 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp 0
transform -1 0 10488 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _234_
timestamp 0
transform 1 0 9660 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _235_
timestamp 0
transform -1 0 17756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _236_
timestamp 0
transform -1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 0
transform -1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _238_
timestamp 0
transform -1 0 17296 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _239_
timestamp 0
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _240_
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _241_
timestamp 0
transform 1 0 7912 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 0
transform -1 0 7360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _243_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _244_
timestamp 0
transform -1 0 8464 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _245_
timestamp 0
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _246_
timestamp 0
transform -1 0 8740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _247_
timestamp 0
transform -1 0 8556 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _248_
timestamp 0
transform 1 0 17388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _249_
timestamp 0
transform -1 0 17112 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _250_
timestamp 0
transform 1 0 17112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _251_
timestamp 0
transform -1 0 16928 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _252_
timestamp 0
transform 1 0 9384 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 0
transform -1 0 8832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 0
transform -1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _256_
timestamp 0
transform -1 0 13064 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 0
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 0
transform -1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _259_
timestamp 0
transform 1 0 12052 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _260_
timestamp 0
transform -1 0 13156 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _261_
timestamp 0
transform -1 0 13340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 0
transform -1 0 13616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _263_
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 0
transform 1 0 10028 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _265_
timestamp 0
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 0
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _267_
timestamp 0
transform -1 0 9568 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _268_
timestamp 0
transform -1 0 17940 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _269_
timestamp 0
transform -1 0 17940 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 0
transform 1 0 15732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 0
transform 1 0 16100 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 0
transform 1 0 15732 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _273_
timestamp 0
transform 1 0 16100 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _274_
timestamp 0
transform 1 0 14904 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _275_
timestamp 0
transform -1 0 16008 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _279_
timestamp 0
transform -1 0 16468 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _280_
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _281_
timestamp 0
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 0
transform -1 0 15916 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 0
transform -1 0 17940 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 0
transform 1 0 11776 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _285_
timestamp 0
transform -1 0 10212 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _286_
timestamp 0
transform 1 0 8372 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _287_
timestamp 0
transform 1 0 10212 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _288_
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _289_
timestamp 0
transform -1 0 14628 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _290_
timestamp 0
transform -1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _291_
timestamp 0
transform 1 0 6992 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _292_
timestamp 0
transform 1 0 8188 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _293_
timestamp 0
transform 1 0 8924 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _294_
timestamp 0
transform 1 0 9384 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _296_
timestamp 0
transform 1 0 11776 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _297_
timestamp 0
transform -1 0 13984 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _298_
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _299_
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _300_
timestamp 0
transform 1 0 11684 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _301_
timestamp 0
transform -1 0 14168 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _302_
timestamp 0
transform 1 0 9384 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _303_
timestamp 0
transform 1 0 7544 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 0
transform -1 0 9384 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _305_
timestamp 0
transform -1 0 6256 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp 0
transform 1 0 6072 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp 0
transform 1 0 5244 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _308_
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _309_
timestamp 0
transform 1 0 7176 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _310_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _311_
timestamp 0
transform -1 0 6808 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _312_
timestamp 0
transform 1 0 3220 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _313_
timestamp 0
transform -1 0 8188 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _314_
timestamp 0
transform 1 0 3864 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 0
transform 1 0 6532 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 0
transform -1 0 7176 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _318_
timestamp 0
transform 1 0 4048 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 0
transform -1 0 3220 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 0
transform -1 0 4600 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 0
transform 1 0 3772 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 0
transform 1 0 3680 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 0
transform -1 0 5612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _329_
timestamp 0
transform 1 0 1932 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _330_
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _331_
timestamp 0
transform -1 0 3220 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 11408 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 0
transform -1 0 6072 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 0
transform -1 0 8832 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 0
transform -1 0 6440 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 0
transform -1 0 8832 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 0
transform -1 0 13984 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 0
transform 1 0 14628 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 0
transform -1 0 13616 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 0
transform 1 0 15916 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_1  clkload0
timestamp 0
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  clkload1
timestamp 0
transform 1 0 4324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp 0
transform 1 0 12512 0 -1 7616
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload3
timestamp 0
transform 1 0 14260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__bufinv_16  clkload4
timestamp 0
transform 1 0 11776 0 -1 15232
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload5
timestamp 0
transform 1 0 14904 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 0
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_162
timestamp 0
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_74
timestamp 0
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 0
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_101
timestamp 0
transform 1 0 10396 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_113
timestamp 0
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_125
timestamp 0
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 0
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_149
timestamp 0
transform 1 0 14812 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_173
timestamp 0
transform 1 0 17020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_181
timestamp 0
transform 1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_34
timestamp 0
transform 1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_65
timestamp 0
transform 1 0 7084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 0
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_120
timestamp 0
transform 1 0 12144 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_178
timestamp 0
transform 1 0 17480 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_182
timestamp 0
transform 1 0 17848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_35
timestamp 0
transform 1 0 4324 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_50
timestamp 0
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_58
timestamp 0
transform 1 0 6440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_64
timestamp 0
transform 1 0 6992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 0
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_92
timestamp 0
transform 1 0 9568 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_114
timestamp 0
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_118
timestamp 0
transform 1 0 11960 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_126
timestamp 0
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 0
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_171
timestamp 0
transform 1 0 16836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_29
timestamp 0
transform 1 0 3772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_41
timestamp 0
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 0
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 0
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_126
timestamp 0
transform 1 0 12696 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_134
timestamp 0
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_157
timestamp 0
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 0
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_11
timestamp 0
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_93
timestamp 0
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_151
timestamp 0
transform 1 0 14996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_103
timestamp 0
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_121
timestamp 0
transform 1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_154
timestamp 0
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 0
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_176
timestamp 0
transform 1 0 17296 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_182
timestamp 0
transform 1 0 17848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_17
timestamp 0
transform 1 0 2668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 0
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_39
timestamp 0
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_43
timestamp 0
transform 1 0 5060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_117
timestamp 0
transform 1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_148
timestamp 0
transform 1 0 14720 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_156
timestamp 0
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_179
timestamp 0
transform 1 0 17572 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_21
timestamp 0
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 0
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 0
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 0
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_121
timestamp 0
transform 1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_130
timestamp 0
transform 1 0 13064 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_142
timestamp 0
transform 1 0 14168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_172
timestamp 0
transform 1 0 16928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_180
timestamp 0
transform 1 0 17664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_23
timestamp 0
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp 0
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_111
timestamp 0
transform 1 0 11316 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_119
timestamp 0
transform 1 0 12052 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_161
timestamp 0
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_11
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_17
timestamp 0
transform 1 0 2668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_25
timestamp 0
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_48
timestamp 0
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_64
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_86
timestamp 0
transform 1 0 9016 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_94
timestamp 0
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_100
timestamp 0
transform 1 0 10304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_133
timestamp 0
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_145
timestamp 0
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_157
timestamp 0
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 0
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 0
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_44
timestamp 0
transform 1 0 5152 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_52
timestamp 0
transform 1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_67
timestamp 0
transform 1 0 7268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 0
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_106
timestamp 0
transform 1 0 10856 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_118
timestamp 0
transform 1 0 11960 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_128
timestamp 0
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_161
timestamp 0
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_23
timestamp 0
transform 1 0 3220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 0
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_63
timestamp 0
transform 1 0 6900 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_75
timestamp 0
transform 1 0 8004 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_87
timestamp 0
transform 1 0 9108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_95
timestamp 0
transform 1 0 9844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_104
timestamp 0
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_143
timestamp 0
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_162
timestamp 0
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_175
timestamp 0
transform 1 0 17204 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_9
timestamp 0
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_62
timestamp 0
transform 1 0 6808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 0
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_89
timestamp 0
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_113
timestamp 0
transform 1 0 11500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 0
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_150
timestamp 0
transform 1 0 14904 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_162
timestamp 0
transform 1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_172
timestamp 0
transform 1 0 16928 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_180
timestamp 0
transform 1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_11
timestamp 0
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_18
timestamp 0
transform 1 0 2760 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_29
timestamp 0
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_41
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 0
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_89
timestamp 0
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_136
timestamp 0
transform 1 0 13616 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_21
timestamp 0
transform 1 0 3036 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_49
timestamp 0
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_61
timestamp 0
transform 1 0 6716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_73
timestamp 0
transform 1 0 7820 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_131
timestamp 0
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_179
timestamp 0
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 0
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_64
timestamp 0
transform 1 0 6992 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_76
timestamp 0
transform 1 0 8096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_84
timestamp 0
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_117
timestamp 0
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_121
timestamp 0
transform 1 0 12236 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 0
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_17
timestamp 0
transform 1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_25
timestamp 0
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_37
timestamp 0
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_44
timestamp 0
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_56
timestamp 0
transform 1 0 6256 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_92
timestamp 0
transform 1 0 9568 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_161
timestamp 0
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_18
timestamp 0
transform 1 0 2760 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_23
timestamp 0
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_35
timestamp 0
transform 1 0 4324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_77
timestamp 0
transform 1 0 8188 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_89
timestamp 0
transform 1 0 9292 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_101
timestamp 0
transform 1 0 10396 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_107
timestamp 0
transform 1 0 10948 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_121
timestamp 0
transform 1 0 12236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_133
timestamp 0
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_145
timestamp 0
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_156
timestamp 0
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_177
timestamp 0
transform 1 0 17388 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_9
timestamp 0
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_18
timestamp 0
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 0
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_58
timestamp 0
transform 1 0 6440 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_93
timestamp 0
transform 1 0 9660 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_105
timestamp 0
transform 1 0 10764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_113
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 0
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_181
timestamp 0
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_23
timestamp 0
transform 1 0 3220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_29
timestamp 0
transform 1 0 3772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_64
timestamp 0
transform 1 0 6992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_76
timestamp 0
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 0
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_140
timestamp 0
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_162
timestamp 0
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_11
timestamp 0
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_23
timestamp 0
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_48
timestamp 0
transform 1 0 5520 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_52
timestamp 0
transform 1 0 5888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_58
timestamp 0
transform 1 0 6440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 0
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_90
timestamp 0
transform 1 0 9384 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_98
timestamp 0
transform 1 0 10120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 0
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_150
timestamp 0
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_162
timestamp 0
transform 1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_38
timestamp 0
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_50
timestamp 0
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_139
timestamp 0
transform 1 0 13892 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 0
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_42
timestamp 0
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_66
timestamp 0
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_75
timestamp 0
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_100
timestamp 0
transform 1 0 10304 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_112
timestamp 0
transform 1 0 11408 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_128
timestamp 0
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_23
timestamp 0
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_35
timestamp 0
transform 1 0 4324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 0
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_65
timestamp 0
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_74
timestamp 0
transform 1 0 7912 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_78
timestamp 0
transform 1 0 8280 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_99
timestamp 0
transform 1 0 10212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_157
timestamp 0
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 0
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_11
timestamp 0
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_25
timestamp 0
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_37
timestamp 0
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_50
timestamp 0
transform 1 0 5704 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_62
timestamp 0
transform 1 0 6808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_102
timestamp 0
transform 1 0 10488 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_108
timestamp 0
transform 1 0 11040 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_136
timestamp 0
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_161
timestamp 0
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_29
timestamp 0
transform 1 0 3772 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 0
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_77
timestamp 0
transform 1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 0
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_117
timestamp 0
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_139
timestamp 0
transform 1 0 13892 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_164
timestamp 0
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_176
timestamp 0
transform 1 0 17296 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_6
timestamp 0
transform 1 0 1656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_10
timestamp 0
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_23
timestamp 0
transform 1 0 3220 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_34
timestamp 0
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_40
timestamp 0
transform 1 0 4784 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_46
timestamp 0
transform 1 0 5336 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_52
timestamp 0
transform 1 0 5888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_60
timestamp 0
transform 1 0 6624 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_64
timestamp 0
transform 1 0 6992 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_70
timestamp 0
transform 1 0 7544 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_76
timestamp 0
transform 1 0 8096 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 0
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_88
timestamp 0
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_94
timestamp 0
transform 1 0 9752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_100
timestamp 0
transform 1 0 10304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_106
timestamp 0
transform 1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_113
timestamp 0
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_118
timestamp 0
transform 1 0 11960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_124
timestamp 0
transform 1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_130
timestamp 0
transform 1 0 13064 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 0
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_144
timestamp 0
transform 1 0 14352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_148
timestamp 0
transform 1 0 14720 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_154
timestamp 0
transform 1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_160
timestamp 0
transform 1 0 15824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_166
timestamp 0
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_172
timestamp 0
transform 1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_178
timestamp 0
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 6716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 7268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform 1 0 7820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 9476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform 1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform -1 0 11408 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 0
transform -1 0 11960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 0
transform 1 0 1748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 0
transform -1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 0
transform -1 0 13064 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 0
transform -1 0 14720 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 0
transform -1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 0
transform 1 0 15548 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 0
transform -1 0 16376 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 0
transform -1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 0
transform 1 0 17204 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 0
transform 1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 0
transform 1 0 17664 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 0
transform 1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 0
transform -1 0 2852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 0
transform -1 0 3680 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 0
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 0
transform -1 0 4784 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 0
transform -1 0 5336 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 0
transform -1 0 5888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 0
transform -1 0 6624 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input33
timestamp 0
transform 1 0 14536 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  output34
timestamp 0
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 18216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 18216 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 18216 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 18216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 18216 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 18216 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 18216 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 18216 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 18216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 18216 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 18216 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 18216 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 18216 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 18216 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 18216 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 18216 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 18216 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 18216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 18216 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_69
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_70
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_72
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_75
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_79
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_87
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_93
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_96
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_97
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_102
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_103
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_105
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_106
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_108
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_111
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_114
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_117
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_120
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_121
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_123
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_124
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_126
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_127
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_129
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_130
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_132
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_133
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_135
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_136
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_138
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_139
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_141
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_142
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_144
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_145
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_147
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_148
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_151
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_155
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_156
timestamp 0
transform 1 0 6256 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_157
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_158
timestamp 0
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_160
timestamp 0
transform 1 0 16560 0 1 18496
box -38 -48 130 592
<< labels >>
rlabel metal1 s 9660 18496 9660 18496 4 VGND
rlabel metal1 s 9660 19040 9660 19040 4 VPWR
rlabel metal2 s 16790 14280 16790 14280 4 _000_
rlabel metal1 s 17480 10710 17480 10710 4 _001_
rlabel metal2 s 10258 17850 10258 17850 4 _002_
rlabel metal2 s 10442 17850 10442 17850 4 _003_
rlabel metal1 s 10120 16626 10120 16626 4 _004_
rlabel metal2 s 17710 9180 17710 9180 4 _005_
rlabel metal1 s 17020 8806 17020 8806 4 _006_
rlabel metal2 s 16974 7786 16974 7786 4 _007_
rlabel metal1 s 7130 8976 7130 8976 4 _008_
rlabel metal2 s 17066 8840 17066 8840 4 _009_
rlabel metal1 s 7406 8942 7406 8942 4 _010_
rlabel metal1 s 6946 9146 6946 9146 4 _011_
rlabel metal1 s 8464 12206 8464 12206 4 _012_
rlabel metal1 s 8970 11866 8970 11866 4 _013_
rlabel metal1 s 8464 11186 8464 11186 4 _014_
rlabel metal1 s 17388 12954 17388 12954 4 _015_
rlabel metal2 s 17158 13328 17158 13328 4 _016_
rlabel metal1 s 17020 11186 17020 11186 4 _017_
rlabel metal2 s 9430 7004 9430 7004 4 _018_
rlabel metal1 s 8832 6630 8832 6630 4 _019_
rlabel metal1 s 8832 5746 8832 5746 4 _020_
rlabel metal1 s 13892 7378 13892 7378 4 _021_
rlabel metal1 s 13248 6426 13248 6426 4 _022_
rlabel metal1 s 13754 7174 13754 7174 4 _023_
rlabel metal2 s 13386 11594 13386 11594 4 _024_
rlabel metal1 s 13386 11254 13386 11254 4 _025_
rlabel metal1 s 12972 10098 12972 10098 4 _026_
rlabel metal2 s 9338 14994 9338 14994 4 _027_
rlabel metal2 s 9614 14620 9614 14620 4 _028_
rlabel metal2 s 9246 14348 9246 14348 4 _029_
rlabel metal1 s 14306 18394 14306 18394 4 _030_
rlabel metal2 s 13662 15674 13662 15674 4 _031_
rlabel metal2 s 12742 15946 12742 15946 4 _032_
rlabel metal1 s 13340 15538 13340 15538 4 _033_
rlabel metal1 s 7636 17714 7636 17714 4 _034_
rlabel metal1 s 7544 17306 7544 17306 4 _035_
rlabel metal2 s 7682 16796 7682 16796 4 _036_
rlabel metal1 s 12742 18292 12742 18292 4 _037_
rlabel metal1 s 2438 11696 2438 11696 4 _038_
rlabel metal1 s 12926 18190 12926 18190 4 _039_
rlabel metal2 s 12834 17952 12834 17952 4 _040_
rlabel metal2 s 2622 8058 2622 8058 4 _041_
rlabel metal2 s 2346 8636 2346 8636 4 _042_
rlabel metal1 s 2162 7718 2162 7718 4 _043_
rlabel metal1 s 15410 18054 15410 18054 4 _044_
rlabel metal2 s 15686 17646 15686 17646 4 _045_
rlabel metal1 s 16422 18190 16422 18190 4 _046_
rlabel metal2 s 4646 17340 4646 17340 4 _047_
rlabel metal1 s 5336 17170 5336 17170 4 _048_
rlabel metal2 s 4830 16796 4830 16796 4 _049_
rlabel metal1 s 14582 14892 14582 14892 4 _050_
rlabel metal1 s 15364 15130 15364 15130 4 _051_
rlabel metal2 s 14766 15844 14766 15844 4 _052_
rlabel metal1 s 3312 11118 3312 11118 4 _053_
rlabel metal2 s 2714 11322 2714 11322 4 _054_
rlabel metal2 s 3450 11492 3450 11492 4 _055_
rlabel metal1 s 14858 10642 14858 10642 4 _056_
rlabel metal1 s 15364 10778 15364 10778 4 _057_
rlabel metal2 s 14766 11492 14766 11492 4 _058_
rlabel metal1 s 2622 17612 2622 17612 4 _059_
rlabel metal2 s 3082 18156 3082 18156 4 _060_
rlabel metal1 s 3082 17102 3082 17102 4 _061_
rlabel metal2 s 15594 5984 15594 5984 4 _062_
rlabel metal1 s 14858 6766 14858 6766 4 _063_
rlabel metal2 s 15226 7174 15226 7174 4 _064_
rlabel metal1 s 14812 7514 14812 7514 4 _065_
rlabel metal1 s 16974 4624 16974 4624 4 _066_
rlabel metal2 s 16698 5066 16698 5066 4 _067_
rlabel metal1 s 17020 4794 17020 4794 4 _068_
rlabel metal1 s 2484 13906 2484 13906 4 _069_
rlabel metal2 s 4830 14382 4830 14382 4 _070_
rlabel metal1 s 2714 13940 2714 13940 4 _071_
rlabel metal2 s 2530 13532 2530 13532 4 _072_
rlabel metal1 s 3726 6324 3726 6324 4 _073_
rlabel metal2 s 3450 5644 3450 5644 4 _074_
rlabel metal2 s 3910 5610 3910 5610 4 _075_
rlabel metal1 s 4738 9894 4738 9894 4 _076_
rlabel metal1 s 5704 8602 5704 8602 4 _077_
rlabel metal1 s 4738 7922 4738 7922 4 _078_
rlabel metal2 s 12190 13532 12190 13532 4 _079_
rlabel metal2 s 12006 13260 12006 13260 4 _080_
rlabel metal1 s 12282 12954 12282 12954 4 _081_
rlabel metal2 s 10810 8636 10810 8636 4 _082_
rlabel metal2 s 10534 8976 10534 8976 4 _083_
rlabel metal2 s 10442 7786 10442 7786 4 _084_
rlabel metal1 s 6762 5644 6762 5644 4 _085_
rlabel metal1 s 6946 5712 6946 5712 4 _086_
rlabel metal1 s 6118 5746 6118 5746 4 _087_
rlabel metal1 s 5290 12852 5290 12852 4 _088_
rlabel metal2 s 5750 13056 5750 13056 4 _089_
rlabel metal1 s 6210 12750 6210 12750 4 _090_
rlabel metal2 s 11270 5066 11270 5066 4 _091_
rlabel metal2 s 11454 5066 11454 5066 4 _092_
rlabel metal2 s 11362 4964 11362 4964 4 _093_
rlabel metal1 s 17480 16082 17480 16082 4 _094_
rlabel metal1 s 17158 15504 17158 15504 4 _095_
rlabel metal2 s 11270 11594 11270 11594 4 _096_
rlabel metal1 s 10534 10778 10534 10778 4 _097_
rlabel metal1 s 10902 10098 10902 10098 4 _098_
rlabel metal1 s 5704 14790 5704 14790 4 _099_
rlabel metal1 s 5658 15436 5658 15436 4 _100_
rlabel metal2 s 6486 15130 6486 15130 4 _101_
rlabel metal1 s 1288 18734 1288 18734 4 a[0]
rlabel metal1 s 6716 18734 6716 18734 4 a[10]
rlabel metal2 s 7314 19805 7314 19805 4 a[11]
rlabel metal2 s 7866 19805 7866 19805 4 a[12]
rlabel metal2 s 8418 19805 8418 19805 4 a[13]
rlabel metal2 s 8970 19805 8970 19805 4 a[14]
rlabel metal2 s 9522 19805 9522 19805 4 a[15]
rlabel metal2 s 10074 19805 10074 19805 4 a[16]
rlabel metal1 s 10580 18734 10580 18734 4 a[17]
rlabel metal1 s 11224 18734 11224 18734 4 a[18]
rlabel metal1 s 11776 18734 11776 18734 4 a[19]
rlabel metal1 s 1748 18734 1748 18734 4 a[1]
rlabel metal2 s 12190 19798 12190 19798 4 a[20]
rlabel metal1 s 12788 18734 12788 18734 4 a[21]
rlabel metal2 s 13570 19805 13570 19805 4 a[22]
rlabel metal1 s 14076 18734 14076 18734 4 a[23]
rlabel metal2 s 14490 19805 14490 19805 4 a[24]
rlabel metal2 s 15042 19805 15042 19805 4 a[25]
rlabel metal2 s 15594 19805 15594 19805 4 a[26]
rlabel metal2 s 16330 19805 16330 19805 4 a[27]
rlabel metal2 s 16882 19805 16882 19805 4 a[28]
rlabel metal2 s 17250 19805 17250 19805 4 a[29]
rlabel metal2 s 2346 19805 2346 19805 4 a[2]
rlabel metal2 s 17710 19798 17710 19798 4 a[30]
rlabel metal1 s 18078 18258 18078 18258 4 a[31]
rlabel metal2 s 2806 19798 2806 19798 4 a[3]
rlabel metal1 s 3496 18734 3496 18734 4 a[4]
rlabel metal1 s 4048 18734 4048 18734 4 a[5]
rlabel metal2 s 4554 19805 4554 19805 4 a[6]
rlabel metal1 s 5060 18734 5060 18734 4 a[7]
rlabel metal2 s 5658 19805 5658 19805 4 a[8]
rlabel metal1 s 6348 18734 6348 18734 4 a[9]
rlabel metal3 s 17603 10676 17603 10676 4 clk
rlabel metal1 s 13570 14280 13570 14280 4 clknet_0_clk
rlabel metal1 s 1564 5746 1564 5746 4 clknet_3_0__leaf_clk
rlabel metal1 s 9108 9010 9108 9010 4 clknet_3_1__leaf_clk
rlabel metal1 s 1426 18156 1426 18156 4 clknet_3_2__leaf_clk
rlabel metal1 s 8418 18224 8418 18224 4 clknet_3_3__leaf_clk
rlabel metal1 s 13156 6290 13156 6290 4 clknet_3_4__leaf_clk
rlabel metal1 s 16054 6834 16054 6834 4 clknet_3_5__leaf_clk
rlabel metal2 s 11868 13294 11868 13294 4 clknet_3_6__leaf_clk
rlabel metal2 s 17894 17170 17894 17170 4 clknet_3_7__leaf_clk
rlabel metal2 s 16146 16320 16146 16320 4 dsa\[0\].last_carry
rlabel metal1 s 17526 15878 17526 15878 4 dsa\[0\].last_carry_next
rlabel metal2 s 16974 11934 16974 11934 4 dsa\[0\].y_out
rlabel metal2 s 17618 14348 17618 14348 4 dsa\[0\].y_out_next
rlabel metal2 s 13294 16252 13294 16252 4 dsa\[10\].last_carry
rlabel metal1 s 12006 15674 12006 15674 4 dsa\[10\].last_carry_next
rlabel metal1 s 13018 15504 13018 15504 4 dsa\[10\].y_in
rlabel metal2 s 12834 13124 12834 13124 4 dsa\[10\].y_out
rlabel metal1 s 14076 12750 14076 12750 4 dsa\[10\].y_out_next
rlabel metal1 s 11316 13906 11316 13906 4 dsa\[11\].last_carry
rlabel metal1 s 11822 13226 11822 13226 4 dsa\[11\].last_carry_next
rlabel metal2 s 9338 13838 9338 13838 4 dsa\[11\].y_out
rlabel metal1 s 11822 13430 11822 13430 4 dsa\[11\].y_out_next
rlabel metal1 s 10258 14960 10258 14960 4 dsa\[12\].last_carry
rlabel metal2 s 8970 14756 8970 14756 4 dsa\[12\].last_carry_next
rlabel metal1 s 10488 12614 10488 12614 4 dsa\[12\].y_out
rlabel metal2 s 9246 13022 9246 13022 4 dsa\[12\].y_out_next
rlabel metal2 s 10902 11764 10902 11764 4 dsa\[13\].last_carry
rlabel metal1 s 9844 10778 9844 10778 4 dsa\[13\].last_carry_next
rlabel metal1 s 12880 10030 12880 10030 4 dsa\[13\].y_out
rlabel metal2 s 11822 9758 11822 9758 4 dsa\[13\].y_out_next
rlabel metal2 s 13570 12036 13570 12036 4 dsa\[14\].last_carry
rlabel metal1 s 12190 11322 12190 11322 4 dsa\[14\].last_carry_next
rlabel metal2 s 10166 8602 10166 8602 4 dsa\[14\].y_out
rlabel metal2 s 13662 9384 13662 9384 4 dsa\[14\].y_out_next
rlabel metal2 s 10718 9350 10718 9350 4 dsa\[15\].last_carry
rlabel metal1 s 9706 8602 9706 8602 4 dsa\[15\].last_carry_next
rlabel metal2 s 12282 6426 12282 6426 4 dsa\[15\].y_out
rlabel metal2 s 10159 6970 10159 6970 4 dsa\[15\].y_out_next
rlabel metal1 s 13570 6800 13570 6800 4 dsa\[16\].last_carry
rlabel metal2 s 12006 6562 12006 6562 4 dsa\[16\].last_carry_next
rlabel metal1 s 11454 5202 11454 5202 4 dsa\[16\].y_out
rlabel metal2 s 13846 5406 13846 5406 4 dsa\[16\].y_out_next
rlabel metal1 s 10994 5712 10994 5712 4 dsa\[17\].last_carry
rlabel metal1 s 10120 4794 10120 4794 4 dsa\[17\].last_carry_next
rlabel metal2 s 9338 6222 9338 6222 4 dsa\[17\].y_out
rlabel metal1 s 11132 5066 11132 5066 4 dsa\[17\].y_out_next
rlabel metal1 s 8740 6766 8740 6766 4 dsa\[18\].last_carry
rlabel metal1 s 9338 6970 9338 6970 4 dsa\[18\].last_carry_next
rlabel metal2 s 5290 5338 5290 5338 4 dsa\[18\].y_out
rlabel metal1 s 6716 5270 6716 5270 4 dsa\[18\].y_out_next
rlabel metal2 s 7774 5202 7774 5202 4 dsa\[19\].last_carry
rlabel metal2 s 6394 4828 6394 4828 4 dsa\[19\].last_carry_next
rlabel metal1 s 6854 8942 6854 8942 4 dsa\[19\].y_out
rlabel metal2 s 5566 6290 5566 6290 4 dsa\[19\].y_out_next
rlabel metal1 s 17572 12818 17572 12818 4 dsa\[1\].last_carry
rlabel metal2 s 16698 12342 16698 12342 4 dsa\[1\].last_carry_next
rlabel metal2 s 16606 9418 16606 9418 4 dsa\[1\].y_out
rlabel metal2 s 16422 10540 16422 10540 4 dsa\[1\].y_out_next
rlabel metal2 s 7590 8500 7590 8500 4 dsa\[20\].last_carry
rlabel metal1 s 5520 7786 5520 7786 4 dsa\[20\].last_carry_next
rlabel metal1 s 8326 11084 8326 11084 4 dsa\[20\].y_out
rlabel metal1 s 6946 9656 6946 9656 4 dsa\[20\].y_out_next
rlabel metal2 s 8142 12036 8142 12036 4 dsa\[21\].last_carry
rlabel metal1 s 7452 11662 7452 11662 4 dsa\[21\].last_carry_next
rlabel metal1 s 5382 12716 5382 12716 4 dsa\[21\].y_out
rlabel metal1 s 6578 11186 6578 11186 4 dsa\[21\].y_out_next
rlabel metal1 s 5198 12614 5198 12614 4 dsa\[22\].last_carry
rlabel metal1 s 4324 12750 4324 12750 4 dsa\[22\].last_carry_next
rlabel metal1 s 6486 14042 6486 14042 4 dsa\[22\].y_out
rlabel metal1 s 7406 12954 7406 12954 4 dsa\[22\].y_out_next
rlabel metal1 s 5612 15130 5612 15130 4 dsa\[23\].last_carry
rlabel metal1 s 4646 14042 4646 14042 4 dsa\[23\].last_carry_next
rlabel metal1 s 7498 16558 7498 16558 4 dsa\[23\].y_out
rlabel metal2 s 6946 15266 6946 15266 4 dsa\[23\].y_out_next
rlabel metal1 s 7912 17646 7912 17646 4 dsa\[24\].last_carry
rlabel metal2 s 6946 18088 6946 18088 4 dsa\[24\].last_carry_next
rlabel metal1 s 5060 16558 5060 16558 4 dsa\[24\].y_out
rlabel metal1 s 6946 16626 6946 16626 4 dsa\[24\].y_out_next
rlabel metal1 s 5750 17646 5750 17646 4 dsa\[25\].last_carry
rlabel metal1 s 4416 17306 4416 17306 4 dsa\[25\].last_carry_next
rlabel metal2 s 1426 16966 1426 16966 4 dsa\[25\].y_out
rlabel metal1 s 2990 16626 2990 16626 4 dsa\[25\].y_out_next
rlabel metal2 s 3174 18530 3174 18530 4 dsa\[26\].last_carry
rlabel metal1 s 2070 17850 2070 17850 4 dsa\[26\].last_carry_next
rlabel metal2 s 2346 15130 2346 15130 4 dsa\[26\].y_out
rlabel metal2 s 4278 16592 4278 16592 4 dsa\[26\].y_out_next
rlabel metal2 s 3174 14586 3174 14586 4 dsa\[27\].last_carry
rlabel metal1 s 1886 14586 1886 14586 4 dsa\[27\].last_carry_next
rlabel metal1 s 2254 11118 2254 11118 4 dsa\[27\].y_out
rlabel metal2 s 1702 13022 1702 13022 4 dsa\[27\].y_out_next
rlabel metal2 s 3082 11424 3082 11424 4 dsa\[28\].last_carry
rlabel metal2 s 1702 10846 1702 10846 4 dsa\[28\].last_carry_next
rlabel metal1 s 4508 8398 4508 8398 4 dsa\[28\].y_out
rlabel metal1 s 3910 10710 3910 10710 4 dsa\[28\].y_out_next
rlabel metal1 s 5198 9690 5198 9690 4 dsa\[29\].last_carry
rlabel metal1 s 4094 8602 4094 8602 4 dsa\[29\].last_carry_next
rlabel metal2 s 1978 7514 1978 7514 4 dsa\[29\].y_out
rlabel metal2 s 5290 7582 5290 7582 4 dsa\[29\].y_out_next
rlabel metal1 s 17434 8874 17434 8874 4 dsa\[2\].last_carry
rlabel metal2 s 16054 8364 16054 8364 4 dsa\[2\].last_carry_next
rlabel metal2 s 17250 5916 17250 5916 4 dsa\[2\].y_out
rlabel metal2 s 16790 7072 16790 7072 4 dsa\[2\].y_out_next
rlabel metal1 s 2714 8500 2714 8500 4 dsa\[30\].last_carry
rlabel metal2 s 1702 8466 1702 8466 4 dsa\[30\].last_carry_next
rlabel metal1 s 3220 6290 3220 6290 4 dsa\[30\].y_out
rlabel metal1 s 2208 6902 2208 6902 4 dsa\[30\].y_out_next
rlabel metal2 s 3726 5678 3726 5678 4 dsa\[31\].last_carry
rlabel metal1 s 2162 5746 2162 5746 4 dsa\[31\].last_carry_next
rlabel metal1 s 3634 5100 3634 5100 4 dsa\[31\].y_out_next
rlabel metal1 s 16744 4794 16744 4794 4 dsa\[3\].last_carry
rlabel metal1 s 15272 4522 15272 4522 4 dsa\[3\].last_carry_next
rlabel metal1 s 14490 6834 14490 6834 4 dsa\[3\].y_out
rlabel metal1 s 16721 5066 16721 5066 4 dsa\[3\].y_out_next
rlabel metal2 s 15410 6596 15410 6596 4 dsa\[4\].last_carry
rlabel metal2 s 14030 6494 14030 6494 4 dsa\[4\].last_carry_next
rlabel metal1 s 14904 10574 14904 10574 4 dsa\[4\].y_out
rlabel metal1 s 14306 8058 14306 8058 4 dsa\[4\].y_out_next
rlabel metal2 s 15962 10438 15962 10438 4 dsa\[5\].last_carry
rlabel metal2 s 14398 10268 14398 10268 4 dsa\[5\].last_carry_next
rlabel metal1 s 14904 14994 14904 14994 4 dsa\[5\].y_out
rlabel metal1 s 15456 11866 15456 11866 4 dsa\[5\].y_out_next
rlabel metal2 s 15962 14790 15962 14790 4 dsa\[6\].last_carry
rlabel metal2 s 14398 14552 14398 14552 4 dsa\[6\].last_carry_next
rlabel metal1 s 16146 16762 16146 16762 4 dsa\[6\].y_out
rlabel metal1 s 14398 16490 14398 16490 4 dsa\[6\].y_out_next
rlabel metal1 s 15272 18258 15272 18258 4 dsa\[7\].last_carry
rlabel metal2 s 15502 17442 15502 17442 4 dsa\[7\].last_carry_next
rlabel metal2 s 12282 17850 12282 17850 4 dsa\[7\].y_out
rlabel metal2 s 17618 17850 17618 17850 4 dsa\[7\].y_out_next
rlabel metal2 s 13570 18054 13570 18054 4 dsa\[8\].last_carry
rlabel metal2 s 12098 17884 12098 17884 4 dsa\[8\].last_carry_next
rlabel metal2 s 9798 17476 9798 17476 4 dsa\[8\].y_out
rlabel metal1 s 10534 17238 10534 17238 4 dsa\[8\].y_out_next
rlabel metal1 s 10442 18224 10442 18224 4 dsa\[9\].last_carry
rlabel metal1 s 9108 17850 9108 17850 4 dsa\[9\].last_carry_next
rlabel metal2 s 10534 15912 10534 15912 4 dsa\[9\].y_out_next
rlabel metal1 s 1564 18598 1564 18598 4 net1
rlabel metal1 s 11270 18598 11270 18598 4 net10
rlabel metal1 s 11270 15062 11270 15062 4 net11
rlabel metal1 s 1886 18598 1886 18598 4 net12
rlabel metal1 s 11822 13906 11822 13906 4 net13
rlabel metal2 s 13018 17579 13018 17579 4 net14
rlabel metal2 s 13386 18496 13386 18496 4 net15
rlabel metal2 s 13754 18462 13754 18462 4 net16
rlabel metal1 s 14812 18258 14812 18258 4 net17
rlabel metal1 s 15410 18598 15410 18598 4 net18
rlabel metal1 s 15594 10676 15594 10676 4 net19
rlabel metal1 s 7038 18598 7038 18598 4 net2
rlabel metal1 s 15916 6698 15916 6698 4 net20
rlabel metal2 s 16606 5729 16606 5729 4 net21
rlabel metal1 s 17388 18598 17388 18598 4 net22
rlabel metal1 s 3496 18938 3496 18938 4 net23
rlabel metal1 s 17848 18598 17848 18598 4 net24
rlabel metal1 s 17250 15912 17250 15912 4 net25
rlabel metal1 s 2116 18870 2116 18870 4 net26
rlabel metal2 s 3450 16490 3450 16490 4 net27
rlabel metal2 s 3726 18428 3726 18428 4 net28
rlabel metal1 s 5244 17646 5244 17646 4 net29
rlabel metal1 s 7774 8942 7774 8942 4 net3
rlabel metal1 s 7682 17612 7682 17612 4 net30
rlabel metal1 s 5428 15470 5428 15470 4 net31
rlabel metal1 s 5428 13294 5428 13294 4 net32
rlabel metal2 s 16882 6494 16882 6494 4 net33
rlabel metal1 s 1518 5134 1518 5134 4 net34
rlabel metal2 s 7636 17068 7636 17068 4 net4
rlabel metal1 s 9016 18870 9016 18870 4 net5
rlabel metal1 s 9936 18666 9936 18666 4 net6
rlabel metal2 s 12466 17749 12466 17749 4 net7
rlabel metal2 s 10258 12716 10258 12716 4 net8
rlabel metal1 s 12926 11050 12926 11050 4 net9
rlabel metal2 s 14490 1588 14490 1588 4 rst
rlabel metal3 s 820 15844 820 15844 4 x
rlabel metal3 s 1004 5236 1004 5236 4 y
flabel metal5 s 1056 15716 18264 16116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 9716 18264 10116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3716 18264 4116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 14644 2128 15044 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8644 2128 9044 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2644 2128 3044 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 14976 18264 15376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8976 18264 9376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 2976 18264 3376 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 13904 2128 14304 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7904 2128 8304 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1904 2128 2304 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 1122 20742 1178 21542 0 FreeSans 280 90 0 0 a[0]
port 3 nsew
flabel metal2 s 6642 20742 6698 21542 0 FreeSans 280 90 0 0 a[10]
port 4 nsew
flabel metal2 s 7194 20742 7250 21542 0 FreeSans 280 90 0 0 a[11]
port 5 nsew
flabel metal2 s 7746 20742 7802 21542 0 FreeSans 280 90 0 0 a[12]
port 6 nsew
flabel metal2 s 8298 20742 8354 21542 0 FreeSans 280 90 0 0 a[13]
port 7 nsew
flabel metal2 s 8850 20742 8906 21542 0 FreeSans 280 90 0 0 a[14]
port 8 nsew
flabel metal2 s 9402 20742 9458 21542 0 FreeSans 280 90 0 0 a[15]
port 9 nsew
flabel metal2 s 9954 20742 10010 21542 0 FreeSans 280 90 0 0 a[16]
port 10 nsew
flabel metal2 s 10506 20742 10562 21542 0 FreeSans 280 90 0 0 a[17]
port 11 nsew
flabel metal2 s 11058 20742 11114 21542 0 FreeSans 280 90 0 0 a[18]
port 12 nsew
flabel metal2 s 11610 20742 11666 21542 0 FreeSans 280 90 0 0 a[19]
port 13 nsew
flabel metal2 s 1674 20742 1730 21542 0 FreeSans 280 90 0 0 a[1]
port 14 nsew
flabel metal2 s 12162 20742 12218 21542 0 FreeSans 280 90 0 0 a[20]
port 15 nsew
flabel metal2 s 12714 20742 12770 21542 0 FreeSans 280 90 0 0 a[21]
port 16 nsew
flabel metal2 s 13266 20742 13322 21542 0 FreeSans 280 90 0 0 a[22]
port 17 nsew
flabel metal2 s 13818 20742 13874 21542 0 FreeSans 280 90 0 0 a[23]
port 18 nsew
flabel metal2 s 14370 20742 14426 21542 0 FreeSans 280 90 0 0 a[24]
port 19 nsew
flabel metal2 s 14922 20742 14978 21542 0 FreeSans 280 90 0 0 a[25]
port 20 nsew
flabel metal2 s 15474 20742 15530 21542 0 FreeSans 280 90 0 0 a[26]
port 21 nsew
flabel metal2 s 16026 20742 16082 21542 0 FreeSans 280 90 0 0 a[27]
port 22 nsew
flabel metal2 s 16578 20742 16634 21542 0 FreeSans 280 90 0 0 a[28]
port 23 nsew
flabel metal2 s 17130 20742 17186 21542 0 FreeSans 280 90 0 0 a[29]
port 24 nsew
flabel metal2 s 2226 20742 2282 21542 0 FreeSans 280 90 0 0 a[2]
port 25 nsew
flabel metal2 s 17682 20742 17738 21542 0 FreeSans 280 90 0 0 a[30]
port 26 nsew
flabel metal2 s 18234 20742 18290 21542 0 FreeSans 280 90 0 0 a[31]
port 27 nsew
flabel metal2 s 2778 20742 2834 21542 0 FreeSans 280 90 0 0 a[3]
port 28 nsew
flabel metal2 s 3330 20742 3386 21542 0 FreeSans 280 90 0 0 a[4]
port 29 nsew
flabel metal2 s 3882 20742 3938 21542 0 FreeSans 280 90 0 0 a[5]
port 30 nsew
flabel metal2 s 4434 20742 4490 21542 0 FreeSans 280 90 0 0 a[6]
port 31 nsew
flabel metal2 s 4986 20742 5042 21542 0 FreeSans 280 90 0 0 a[7]
port 32 nsew
flabel metal2 s 5538 20742 5594 21542 0 FreeSans 280 90 0 0 a[8]
port 33 nsew
flabel metal2 s 6090 20742 6146 21542 0 FreeSans 280 90 0 0 a[9]
port 34 nsew
flabel metal3 s 18598 10616 19398 10736 0 FreeSans 600 0 0 0 clk
port 35 nsew
flabel metal2 s 14462 0 14518 800 0 FreeSans 280 90 0 0 rst
port 36 nsew
flabel metal3 s 0 15784 800 15904 0 FreeSans 600 0 0 0 x
port 37 nsew
flabel metal3 s 0 5176 800 5296 0 FreeSans 600 0 0 0 y
port 38 nsew
<< properties >>
string FIXED_BBOX 0 0 19398 21542
<< end >>
